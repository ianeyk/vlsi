magic
tech sky130A
timestamp 1695581597
<< nwell >>
rect -70 445 650 885
<< nmos >>
rect 0 -5 15 395
rect 145 -5 160 395
rect 210 -5 225 395
rect 355 295 370 395
rect 500 295 515 395
rect 565 295 580 395
rect 355 165 370 265
<< pmos >>
rect 0 595 15 695
rect 0 465 15 565
rect 145 465 160 565
rect 210 465 225 565
rect 355 465 370 865
rect 500 465 515 865
rect 565 465 580 865
<< ndiff >>
rect -50 380 0 395
rect -50 10 -35 380
rect -15 10 0 380
rect -50 -5 0 10
rect 15 380 65 395
rect 15 10 30 380
rect 50 10 65 380
rect 15 -5 65 10
rect 95 380 145 395
rect 95 10 110 380
rect 130 10 145 380
rect 95 -5 145 10
rect 160 380 210 395
rect 160 10 175 380
rect 195 10 210 380
rect 160 -5 210 10
rect 225 380 275 395
rect 225 10 240 380
rect 260 10 275 380
rect 305 380 355 395
rect 305 310 320 380
rect 340 310 355 380
rect 305 295 355 310
rect 370 380 420 395
rect 370 310 385 380
rect 405 310 420 380
rect 370 295 420 310
rect 450 380 500 395
rect 450 310 465 380
rect 485 310 500 380
rect 450 295 500 310
rect 515 380 565 395
rect 515 310 530 380
rect 550 310 565 380
rect 515 295 565 310
rect 580 380 630 395
rect 580 310 595 380
rect 615 310 630 380
rect 580 295 630 310
rect 305 250 355 265
rect 305 180 320 250
rect 340 180 355 250
rect 305 165 355 180
rect 370 250 420 265
rect 370 180 385 250
rect 405 180 420 250
rect 370 165 420 180
rect 225 -5 275 10
<< pdiff >>
rect 305 850 355 865
rect -50 680 0 695
rect -50 610 -35 680
rect -15 610 0 680
rect -50 595 0 610
rect 15 680 65 695
rect 15 610 30 680
rect 50 610 65 680
rect 15 595 65 610
rect -50 550 0 565
rect -50 480 -35 550
rect -15 480 0 550
rect -50 465 0 480
rect 15 550 65 565
rect 15 480 30 550
rect 50 480 65 550
rect 15 465 65 480
rect 95 550 145 565
rect 95 480 110 550
rect 130 480 145 550
rect 95 465 145 480
rect 160 550 210 565
rect 160 480 175 550
rect 195 480 210 550
rect 160 465 210 480
rect 225 550 275 565
rect 225 480 240 550
rect 260 480 275 550
rect 225 465 275 480
rect 305 480 320 850
rect 340 480 355 850
rect 305 465 355 480
rect 370 850 420 865
rect 370 480 385 850
rect 405 480 420 850
rect 370 465 420 480
rect 450 850 500 865
rect 450 480 465 850
rect 485 480 500 850
rect 450 465 500 480
rect 515 850 565 865
rect 515 480 530 850
rect 550 480 565 850
rect 515 465 565 480
rect 580 850 630 865
rect 580 480 595 850
rect 615 480 630 850
rect 580 465 630 480
<< ndiffc >>
rect -35 10 -15 380
rect 30 10 50 380
rect 110 10 130 380
rect 175 10 195 380
rect 240 10 260 380
rect 320 310 340 380
rect 385 310 405 380
rect 465 310 485 380
rect 530 310 550 380
rect 595 310 615 380
rect 320 180 340 250
rect 385 180 405 250
<< pdiffc >>
rect -35 610 -15 680
rect 30 610 50 680
rect -35 480 -15 550
rect 30 480 50 550
rect 110 480 130 550
rect 175 480 195 550
rect 240 480 260 550
rect 320 480 340 850
rect 385 480 405 850
rect 465 480 485 850
rect 530 480 550 850
rect 595 480 615 850
<< poly >>
rect 355 865 370 880
rect 500 865 515 880
rect 565 865 580 880
rect 0 695 15 710
rect 185 610 225 620
rect 0 565 15 595
rect 185 590 195 610
rect 215 590 225 610
rect 185 580 225 590
rect 145 565 160 580
rect 210 565 225 580
rect 0 395 15 465
rect 145 450 160 465
rect 210 450 225 465
rect 40 440 185 450
rect 40 420 50 440
rect 70 435 155 440
rect 70 420 80 435
rect 40 410 80 420
rect 145 420 155 435
rect 175 420 185 440
rect 145 410 185 420
rect 210 440 310 450
rect 210 430 280 440
rect 145 395 160 410
rect 210 395 225 430
rect 270 420 280 430
rect 300 420 310 440
rect 270 410 310 420
rect 355 395 370 465
rect 500 450 515 465
rect 395 440 435 450
rect 395 420 405 440
rect 425 425 435 440
rect 500 440 540 450
rect 500 425 510 440
rect 425 420 510 425
rect 530 420 540 440
rect 395 410 540 420
rect 565 425 580 465
rect 625 440 665 450
rect 625 425 635 440
rect 565 420 635 425
rect 655 420 665 440
rect 565 410 665 420
rect 500 395 515 410
rect 565 395 580 410
rect 355 265 370 295
rect 500 280 515 295
rect 565 280 580 295
rect 540 270 580 280
rect 540 250 550 270
rect 570 250 580 270
rect 540 240 580 250
rect 355 150 370 165
rect 355 140 395 150
rect 355 120 365 140
rect 385 120 395 140
rect 355 110 395 120
rect 0 -20 15 -5
rect 145 -20 160 -5
rect 210 -20 225 -5
<< polycont >>
rect 195 590 215 610
rect 50 420 70 440
rect 155 420 175 440
rect 280 420 300 440
rect 405 420 425 440
rect 510 420 530 440
rect 635 420 655 440
rect 550 250 570 270
rect 365 120 385 140
<< locali >>
rect 395 880 540 900
rect 395 860 415 880
rect 520 860 540 880
rect 310 850 350 860
rect -45 680 -5 690
rect -45 610 -35 680
rect -15 610 -5 680
rect -45 600 -5 610
rect 20 680 60 690
rect 20 610 30 680
rect 50 620 60 680
rect 50 610 225 620
rect 20 600 195 610
rect 100 560 120 600
rect 185 590 195 600
rect 215 590 225 610
rect 185 580 225 590
rect -45 550 -5 560
rect -45 480 -35 550
rect -15 480 -5 550
rect -45 470 -5 480
rect 20 550 60 560
rect 20 480 30 550
rect 50 480 60 550
rect 20 470 60 480
rect 40 450 60 470
rect 100 550 140 560
rect 100 480 110 550
rect 130 480 140 550
rect 100 470 140 480
rect 165 550 205 560
rect 165 480 175 550
rect 195 480 205 550
rect 165 470 205 480
rect 230 550 270 560
rect 230 480 240 550
rect 260 480 270 550
rect 230 470 270 480
rect 310 480 320 850
rect 340 480 350 850
rect 310 470 350 480
rect 375 850 415 860
rect 375 480 385 850
rect 405 480 415 850
rect 375 470 415 480
rect 455 850 495 860
rect 455 480 465 850
rect 485 480 495 850
rect 455 470 495 480
rect 520 850 560 860
rect 520 480 530 850
rect 550 480 560 850
rect 520 470 560 480
rect 585 850 625 860
rect 585 480 595 850
rect 615 620 625 850
rect 615 600 665 620
rect 615 480 625 600
rect 585 470 625 480
rect 40 440 80 450
rect 40 420 50 440
rect 70 420 80 440
rect 40 410 80 420
rect 100 390 120 470
rect 230 450 250 470
rect 145 440 250 450
rect 145 420 155 440
rect 175 430 250 440
rect 175 420 185 430
rect 145 410 185 420
rect 230 390 250 430
rect 270 440 310 450
rect 270 420 280 440
rect 300 420 310 440
rect 270 410 310 420
rect 290 390 310 410
rect 395 440 435 450
rect 395 420 405 440
rect 425 420 435 440
rect 395 410 435 420
rect 395 390 415 410
rect -45 380 -5 390
rect -45 10 -35 380
rect -15 10 -5 380
rect -45 0 -5 10
rect 20 380 60 390
rect 20 10 30 380
rect 50 10 60 380
rect 20 0 60 10
rect 100 380 140 390
rect 100 10 110 380
rect 130 10 140 380
rect 100 0 140 10
rect 165 380 205 390
rect 165 10 175 380
rect 195 10 205 380
rect 165 0 205 10
rect 230 380 270 390
rect 230 10 240 380
rect 260 260 270 380
rect 290 380 350 390
rect 290 370 320 380
rect 310 310 320 370
rect 340 310 350 380
rect 310 300 350 310
rect 375 380 415 390
rect 375 310 385 380
rect 405 310 415 380
rect 375 300 415 310
rect 455 390 475 470
rect 500 440 540 450
rect 500 420 510 440
rect 530 430 540 440
rect 585 430 605 470
rect 645 450 665 490
rect 530 420 605 430
rect 500 410 605 420
rect 625 440 665 450
rect 625 420 635 440
rect 655 420 665 440
rect 625 410 665 420
rect 585 390 605 410
rect 455 380 495 390
rect 455 310 465 380
rect 485 310 495 380
rect 455 300 495 310
rect 520 380 560 390
rect 520 310 530 380
rect 550 310 560 380
rect 520 300 560 310
rect 585 380 625 390
rect 585 310 595 380
rect 615 310 625 380
rect 585 300 625 310
rect 455 260 475 300
rect 540 270 580 280
rect 540 260 550 270
rect 260 250 350 260
rect 260 240 320 250
rect 260 10 270 240
rect 310 180 320 240
rect 340 180 350 250
rect 310 170 350 180
rect 375 250 550 260
rect 570 250 580 270
rect 375 180 385 250
rect 405 240 580 250
rect 405 180 415 240
rect 375 170 415 180
rect 230 0 270 10
rect 355 140 395 150
rect 355 120 365 140
rect 385 120 395 140
rect 355 110 395 120
rect 40 -20 60 0
rect 165 -20 185 0
rect 40 -40 185 -20
rect 355 -30 375 110
rect 345 -40 385 -30
rect 345 -60 355 -40
rect 375 -60 385 -40
rect 345 -70 385 -60
<< viali >>
rect 175 480 195 550
rect 320 480 340 850
rect -35 10 -15 380
rect 530 310 550 380
rect 355 -60 375 -40
<< metal1 >>
rect -50 850 665 860
rect -50 550 320 850
rect -50 480 175 550
rect 195 480 320 550
rect 340 480 665 850
rect -50 470 665 480
rect -50 380 665 390
rect -50 10 -35 380
rect -15 310 530 380
rect 550 310 665 380
rect -15 10 665 310
rect -50 0 665 10
rect -50 -40 665 -30
rect -50 -45 355 -40
rect 345 -60 355 -45
rect 375 -45 665 -40
rect 375 -60 385 -45
rect 345 -70 385 -60
<< end >>
