magic
tech sky130A
timestamp 1697171622
<< nwell >>
rect 2895 880 3115 1570
rect 3020 875 3115 880
<< locali >>
rect 2905 2415 3060 2435
rect 2905 960 2925 2415
rect 2970 2145 3060 2155
rect 2970 2125 2980 2145
rect 3000 2135 3060 2145
rect 3000 2125 3010 2135
rect 2970 2115 3010 2125
rect 2970 1700 3010 1710
rect 2970 1680 2980 1700
rect 3000 1690 3010 1700
rect 3000 1680 3060 1690
rect 2970 1670 3060 1680
rect 2965 1595 3060 1615
rect 2965 1030 2985 1595
rect 2945 1020 2985 1030
rect 2945 1000 2955 1020
rect 2975 1000 2985 1020
rect 2945 990 2985 1000
rect 3005 1190 3060 1210
rect 2905 950 2985 960
rect 2905 940 2955 950
rect 2945 930 2955 940
rect 2975 930 2985 950
rect 2945 920 2985 930
rect 3005 900 3025 1190
rect 2855 880 3025 900
rect 2855 790 3025 810
rect 3005 375 3025 790
rect 3005 355 3060 375
<< viali >>
rect 2980 2125 3000 2145
rect 2980 1680 3000 1700
rect 2955 1000 2975 1020
rect 2955 930 2975 950
<< metal1 >>
rect 2970 2145 3010 2155
rect 2970 2125 2980 2145
rect 3000 2125 3010 2145
rect 2970 2115 3010 2125
rect 3040 1755 3055 2340
rect 2970 1700 3010 1710
rect 2970 1680 2980 1700
rect 3000 1680 3010 1700
rect 2970 1670 3010 1680
rect 2860 1550 2875 1650
rect 2860 1250 3055 1550
rect 2860 900 2875 1250
rect 2945 1020 2985 1030
rect 2945 1005 2955 1020
rect 2905 1000 2955 1005
rect 2975 1000 2985 1020
rect 2905 990 2985 1000
rect 2905 865 2920 990
rect 2855 850 2920 865
rect 2945 950 2985 960
rect 2945 930 2955 950
rect 2975 930 2985 950
rect 2945 920 2985 930
rect 2945 835 2960 920
rect 2855 820 2960 835
rect 2860 340 2875 790
rect 2860 40 3055 340
use bias  bias_0
timestamp 1697165931
transform 1 0 785 0 1 80
box -780 -75 2110 1605
use opamp  opamp_0
timestamp 1697128104
transform 1 0 3090 0 1 410
box -70 -435 1410 2025
<< labels >>
flabel metal1 2970 1690 2970 1690 7 FreeSans 160 0 0 0 V1
port 1 w
flabel metal1 2970 2135 2970 2135 7 FreeSans 160 0 0 0 V2
port 2 w
flabel space 4500 600 4500 600 3 FreeSans 160 0 0 0 Vout
port 3 e
flabel space 25 875 25 875 7 FreeSans 160 0 0 0 Ib
port 4 w
flabel space 25 1255 25 1255 7 FreeSans 160 0 0 0 VP
port 5 w
flabel space 25 435 25 435 7 FreeSans 160 0 0 0 VN
port 6 w
<< end >>
