magic
tech sky130A
timestamp 1694271401
<< nwell >>
rect -120 235 200 475
<< nmos >>
rect -10 0 5 200
rect 55 0 70 200
<< pmos >>
rect 0 255 15 455
rect 65 255 80 455
<< ndiff >>
rect -60 185 -10 200
rect -60 15 -45 185
rect -25 15 -10 185
rect -60 0 -10 15
rect 5 0 55 200
rect 70 185 120 200
rect 70 15 85 185
rect 105 15 120 185
rect 70 0 120 15
<< pdiff >>
rect -50 440 0 455
rect -50 270 -35 440
rect -15 270 0 440
rect -50 255 0 270
rect 15 440 65 455
rect 15 270 30 440
rect 50 270 65 440
rect 15 255 65 270
rect 80 440 130 455
rect 80 270 95 440
rect 115 270 130 440
rect 80 255 130 270
<< ndiffc >>
rect -45 15 -25 185
rect 85 15 105 185
<< pdiffc >>
rect -35 270 -15 440
rect 30 270 50 440
rect 95 270 115 440
<< psubdiff >>
rect -110 185 -60 200
rect -110 15 -95 185
rect -75 15 -60 185
rect -110 0 -60 15
rect 150 185 200 200
rect 150 15 165 185
rect 185 15 200 185
rect 150 0 200 15
<< nsubdiff >>
rect -100 440 -50 455
rect -100 270 -85 440
rect -65 270 -50 440
rect -100 255 -50 270
rect 130 440 180 455
rect 130 270 145 440
rect 165 270 180 440
rect 130 255 180 270
<< psubdiffcont >>
rect -95 15 -75 185
rect 165 15 185 185
<< nsubdiffcont >>
rect -85 270 -65 440
rect 145 270 165 440
<< poly >>
rect 0 455 15 470
rect 65 455 80 470
rect 0 230 15 255
rect 65 230 80 255
rect -10 215 15 230
rect 55 215 80 230
rect -10 200 5 215
rect 55 200 70 215
rect -10 -15 5 0
rect 55 -15 70 0
rect -35 -25 5 -15
rect -35 -45 -25 -25
rect -5 -45 5 -25
rect -35 -55 5 -45
rect 30 -25 70 -15
rect 30 -45 40 -25
rect 60 -45 70 -25
rect 30 -55 70 -45
<< polycont >>
rect -25 -45 -5 -25
rect 40 -45 60 -25
<< locali >>
rect -95 440 -5 450
rect -95 270 -85 440
rect -65 270 -35 440
rect -15 270 -5 440
rect -95 260 -5 270
rect 20 440 60 450
rect 20 270 30 440
rect 50 270 60 440
rect 20 260 60 270
rect 85 440 175 450
rect 85 270 95 440
rect 115 270 145 440
rect 165 270 175 440
rect 85 260 175 270
rect 40 195 60 260
rect -105 185 -15 195
rect -105 15 -95 185
rect -75 15 -45 185
rect -25 15 -15 185
rect 40 185 115 195
rect 40 175 85 185
rect -105 5 -15 15
rect 75 15 85 175
rect 105 15 115 185
rect 75 5 115 15
rect 155 185 195 195
rect 155 15 165 185
rect 185 15 195 185
rect 155 5 195 15
rect 95 -15 115 5
rect -120 -25 5 -15
rect -120 -35 -25 -25
rect -35 -45 -25 -35
rect -5 -45 5 -25
rect -35 -55 5 -45
rect 30 -25 70 -15
rect 30 -45 40 -25
rect 60 -45 70 -25
rect 95 -35 200 -15
rect 30 -55 70 -45
rect 30 -75 50 -55
rect -120 -95 50 -75
<< viali >>
rect -85 270 -65 440
rect -35 270 -15 440
rect 95 270 115 440
rect 145 270 165 440
rect -95 15 -75 185
rect -45 15 -25 185
rect 165 15 185 185
<< metal1 >>
rect -120 440 200 455
rect -120 270 -85 440
rect -65 270 -35 440
rect -15 270 95 440
rect 115 270 145 440
rect 165 270 200 440
rect -120 255 200 270
rect -120 185 200 200
rect -120 15 -95 185
rect -75 15 -45 185
rect -25 15 165 185
rect 185 15 200 185
rect -120 0 200 15
<< labels >>
rlabel locali -120 -25 -120 -25 7 A
port 1 w
rlabel locali -120 -85 -120 -85 7 B
port 2 w
rlabel locali 200 -25 200 -25 3 Y
port 3 e
rlabel metal1 -120 355 -120 355 7 VP
port 4 w
rlabel metal1 -120 100 -120 100 7 VN
port 5 w
<< end >>
