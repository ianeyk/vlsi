magic
tech sky130A
timestamp 1697030486
<< error_p >>
rect 125 2047 145 2050
rect 125 1783 128 2047
rect 142 1783 145 2047
rect 125 1780 145 1783
rect 325 2047 345 2050
rect 325 1783 328 2047
rect 342 1783 345 2047
rect 325 1780 345 1783
rect 525 2047 545 2050
rect 525 1783 528 2047
rect 542 1783 545 2047
rect 525 1780 545 1783
rect 725 2047 745 2050
rect 725 1783 728 2047
rect 742 1783 745 2047
rect 725 1780 745 1783
rect 925 2047 945 2050
rect 925 1783 928 2047
rect 942 1783 945 2047
rect 925 1780 945 1783
rect 1125 2047 1145 2050
rect 1125 1783 1128 2047
rect 1142 1783 1145 2047
rect 1125 1780 1145 1783
rect 125 1577 145 1580
rect 125 1313 128 1577
rect 142 1313 145 1577
rect 125 1310 145 1313
rect 1125 1577 1145 1580
rect 1125 1313 1128 1577
rect 1142 1313 1145 1577
rect 1125 1310 1145 1313
rect 125 1097 145 1100
rect 125 833 128 1097
rect 142 833 145 1097
rect 125 830 145 833
rect 325 1097 345 1100
rect 325 833 328 1097
rect 342 833 345 1097
rect 325 830 345 833
rect 525 1097 545 1100
rect 525 833 528 1097
rect 542 833 545 1097
rect 525 830 545 833
rect 725 1097 745 1100
rect 725 833 728 1097
rect 742 833 745 1097
rect 725 830 745 833
rect 925 1097 945 1100
rect 925 833 928 1097
rect 942 833 945 1097
rect 925 830 945 833
rect 1125 1097 1145 1100
rect 1125 833 1128 1097
rect 1142 833 1145 1097
rect 1125 830 1145 833
rect 125 -123 145 -120
rect 125 -387 128 -123
rect 142 -387 145 -123
rect 125 -390 145 -387
rect 325 -123 345 -120
rect 325 -387 328 -123
rect 342 -387 345 -123
rect 325 -390 345 -387
rect 525 -123 545 -120
rect 525 -387 528 -123
rect 542 -387 545 -123
rect 525 -390 545 -387
rect 725 -123 745 -120
rect 725 -387 728 -123
rect 742 -387 745 -123
rect 725 -390 745 -387
rect 925 -123 945 -120
rect 925 -387 928 -123
rect 942 -387 945 -123
rect 925 -390 945 -387
rect 1125 -123 1145 -120
rect 1125 -387 1128 -123
rect 1142 -387 1145 -123
rect 1125 -390 1145 -387
<< nwell >>
rect 90 780 1180 1135
rect 10 775 1340 780
rect -70 375 1340 775
<< nmos >>
rect 160 1765 210 2065
rect 260 1765 310 2065
rect 360 1765 410 2065
rect 460 1765 510 2065
rect 560 1765 610 2065
rect 660 1765 710 2065
rect 760 1765 810 2065
rect 860 1765 910 2065
rect 960 1765 1010 2065
rect 1060 1765 1110 2065
rect 160 1295 210 1595
rect 260 1295 310 1595
rect 360 1295 410 1595
rect 460 1295 510 1595
rect 560 1295 610 1595
rect 660 1295 710 1595
rect 760 1295 810 1595
rect 860 1295 910 1595
rect 960 1295 1010 1595
rect 1060 1295 1110 1595
rect 0 0 50 300
rect 100 0 150 300
rect 280 0 330 300
rect 380 0 430 300
rect 560 0 610 300
rect 660 0 710 300
rect 840 0 890 300
rect 940 0 990 300
rect 1120 0 1170 300
rect 1220 0 1270 300
rect 160 -405 210 -105
rect 260 -405 310 -105
rect 360 -405 410 -105
rect 460 -405 510 -105
rect 560 -405 610 -105
rect 660 -405 710 -105
rect 760 -405 810 -105
rect 860 -405 910 -105
rect 960 -405 1010 -105
rect 1060 -405 1110 -105
<< pmos >>
rect 160 815 210 1115
rect 260 815 310 1115
rect 360 815 410 1115
rect 460 815 510 1115
rect 560 815 610 1115
rect 660 815 710 1115
rect 760 815 810 1115
rect 860 815 910 1115
rect 960 815 1010 1115
rect 1060 815 1110 1115
rect 0 395 50 695
rect 100 395 150 695
rect 280 395 330 695
rect 380 395 430 695
rect 560 395 610 695
rect 660 395 710 695
rect 840 395 890 695
rect 940 395 990 695
rect 1120 395 1170 695
rect 1220 395 1270 695
<< ndiff >>
rect 110 2050 160 2065
rect 110 1780 125 2050
rect 145 1780 160 2050
rect 110 1765 160 1780
rect 210 2050 260 2065
rect 210 1780 225 2050
rect 245 1780 260 2050
rect 210 1765 260 1780
rect 310 2050 360 2065
rect 310 1780 325 2050
rect 345 1780 360 2050
rect 310 1765 360 1780
rect 410 2050 460 2065
rect 410 1780 425 2050
rect 445 1780 460 2050
rect 410 1765 460 1780
rect 510 2050 560 2065
rect 510 1780 525 2050
rect 545 1780 560 2050
rect 510 1765 560 1780
rect 610 2050 660 2065
rect 610 1780 625 2050
rect 645 1780 660 2050
rect 610 1765 660 1780
rect 710 2050 760 2065
rect 710 1780 725 2050
rect 745 1780 760 2050
rect 710 1765 760 1780
rect 810 2050 860 2065
rect 810 1780 825 2050
rect 845 1780 860 2050
rect 810 1765 860 1780
rect 910 2050 960 2065
rect 910 1780 925 2050
rect 945 1780 960 2050
rect 910 1765 960 1780
rect 1010 2050 1060 2065
rect 1010 1780 1025 2050
rect 1045 1780 1060 2050
rect 1010 1765 1060 1780
rect 1110 2050 1160 2065
rect 1110 1780 1125 2050
rect 1145 1780 1160 2050
rect 1110 1765 1160 1780
rect 110 1580 160 1595
rect 110 1310 125 1580
rect 145 1310 160 1580
rect 110 1295 160 1310
rect 210 1580 260 1595
rect 210 1310 225 1580
rect 245 1310 260 1580
rect 210 1295 260 1310
rect 310 1580 360 1595
rect 310 1310 325 1580
rect 345 1310 360 1580
rect 310 1295 360 1310
rect 410 1580 460 1595
rect 410 1310 425 1580
rect 445 1310 460 1580
rect 410 1295 460 1310
rect 510 1580 560 1595
rect 510 1310 525 1580
rect 545 1310 560 1580
rect 510 1295 560 1310
rect 610 1580 660 1595
rect 610 1310 625 1580
rect 645 1310 660 1580
rect 610 1295 660 1310
rect 710 1580 760 1595
rect 710 1310 725 1580
rect 745 1310 760 1580
rect 710 1295 760 1310
rect 810 1580 860 1595
rect 810 1310 825 1580
rect 845 1310 860 1580
rect 810 1295 860 1310
rect 910 1580 960 1595
rect 910 1310 925 1580
rect 945 1310 960 1580
rect 910 1295 960 1310
rect 1010 1580 1060 1595
rect 1010 1310 1025 1580
rect 1045 1310 1060 1580
rect 1010 1295 1060 1310
rect 1110 1580 1160 1595
rect 1110 1310 1125 1580
rect 1145 1310 1160 1580
rect 1110 1295 1160 1310
rect -50 285 0 300
rect -50 15 -35 285
rect -15 15 0 285
rect -50 0 0 15
rect 50 285 100 300
rect 50 15 65 285
rect 85 15 100 285
rect 50 0 100 15
rect 150 285 200 300
rect 150 15 165 285
rect 185 15 200 285
rect 150 0 200 15
rect 230 285 280 300
rect 230 15 245 285
rect 265 15 280 285
rect 230 0 280 15
rect 330 285 380 300
rect 330 15 345 285
rect 365 15 380 285
rect 330 0 380 15
rect 430 285 480 300
rect 430 15 445 285
rect 465 15 480 285
rect 430 0 480 15
rect 510 285 560 300
rect 510 15 525 285
rect 545 15 560 285
rect 510 0 560 15
rect 610 285 660 300
rect 610 15 625 285
rect 645 15 660 285
rect 610 0 660 15
rect 710 285 760 300
rect 710 15 725 285
rect 745 15 760 285
rect 710 0 760 15
rect 790 285 840 300
rect 790 15 805 285
rect 825 15 840 285
rect 790 0 840 15
rect 890 285 940 300
rect 890 15 905 285
rect 925 15 940 285
rect 890 0 940 15
rect 990 285 1040 300
rect 990 15 1005 285
rect 1025 15 1040 285
rect 990 0 1040 15
rect 1070 285 1120 300
rect 1070 15 1085 285
rect 1105 15 1120 285
rect 1070 0 1120 15
rect 1170 285 1220 300
rect 1170 15 1185 285
rect 1205 15 1220 285
rect 1170 0 1220 15
rect 1270 285 1320 300
rect 1270 15 1285 285
rect 1305 15 1320 285
rect 1270 0 1320 15
rect 110 -120 160 -105
rect 110 -390 125 -120
rect 145 -390 160 -120
rect 110 -405 160 -390
rect 210 -120 260 -105
rect 210 -390 225 -120
rect 245 -390 260 -120
rect 210 -405 260 -390
rect 310 -120 360 -105
rect 310 -390 325 -120
rect 345 -390 360 -120
rect 310 -405 360 -390
rect 410 -120 460 -105
rect 410 -390 425 -120
rect 445 -390 460 -120
rect 410 -405 460 -390
rect 510 -120 560 -105
rect 510 -390 525 -120
rect 545 -390 560 -120
rect 510 -405 560 -390
rect 610 -120 660 -105
rect 610 -390 625 -120
rect 645 -390 660 -120
rect 610 -405 660 -390
rect 710 -120 760 -105
rect 710 -390 725 -120
rect 745 -390 760 -120
rect 710 -405 760 -390
rect 810 -120 860 -105
rect 810 -390 825 -120
rect 845 -390 860 -120
rect 810 -405 860 -390
rect 910 -120 960 -105
rect 910 -390 925 -120
rect 945 -390 960 -120
rect 910 -405 960 -390
rect 1010 -120 1060 -105
rect 1010 -390 1025 -120
rect 1045 -390 1060 -120
rect 1010 -405 1060 -390
rect 1110 -120 1160 -105
rect 1110 -390 1125 -120
rect 1145 -390 1160 -120
rect 1110 -405 1160 -390
<< pdiff >>
rect 110 1100 160 1115
rect 110 830 125 1100
rect 145 830 160 1100
rect 110 815 160 830
rect 210 1100 260 1115
rect 210 830 225 1100
rect 245 830 260 1100
rect 210 815 260 830
rect 310 1100 360 1115
rect 310 830 325 1100
rect 345 830 360 1100
rect 310 815 360 830
rect 410 1100 460 1115
rect 410 830 425 1100
rect 445 830 460 1100
rect 410 815 460 830
rect 510 1100 560 1115
rect 510 830 525 1100
rect 545 830 560 1100
rect 510 815 560 830
rect 610 1100 660 1115
rect 610 830 625 1100
rect 645 830 660 1100
rect 610 815 660 830
rect 710 1100 760 1115
rect 710 830 725 1100
rect 745 830 760 1100
rect 710 815 760 830
rect 810 1100 860 1115
rect 810 830 825 1100
rect 845 830 860 1100
rect 810 815 860 830
rect 910 1100 960 1115
rect 910 830 925 1100
rect 945 830 960 1100
rect 910 815 960 830
rect 1010 1100 1060 1115
rect 1010 830 1025 1100
rect 1045 830 1060 1100
rect 1010 815 1060 830
rect 1110 1100 1160 1115
rect 1110 830 1125 1100
rect 1145 830 1160 1100
rect 1110 815 1160 830
rect -50 680 0 695
rect -50 410 -35 680
rect -15 410 0 680
rect -50 395 0 410
rect 50 680 100 695
rect 50 410 65 680
rect 85 410 100 680
rect 50 395 100 410
rect 150 680 200 695
rect 150 410 165 680
rect 185 410 200 680
rect 150 395 200 410
rect 230 680 280 695
rect 230 410 245 680
rect 265 410 280 680
rect 230 395 280 410
rect 330 680 380 695
rect 330 410 345 680
rect 365 410 380 680
rect 330 395 380 410
rect 430 680 480 695
rect 430 410 445 680
rect 465 410 480 680
rect 430 395 480 410
rect 510 680 560 695
rect 510 410 525 680
rect 545 410 560 680
rect 510 395 560 410
rect 610 680 660 695
rect 610 410 625 680
rect 645 410 660 680
rect 610 395 660 410
rect 710 680 760 695
rect 710 410 725 680
rect 745 410 760 680
rect 710 395 760 410
rect 790 680 840 695
rect 790 410 805 680
rect 825 410 840 680
rect 790 395 840 410
rect 890 680 940 695
rect 890 410 905 680
rect 925 410 940 680
rect 890 395 940 410
rect 990 680 1040 695
rect 990 410 1005 680
rect 1025 410 1040 680
rect 990 395 1040 410
rect 1070 680 1120 695
rect 1070 410 1085 680
rect 1105 410 1120 680
rect 1070 395 1120 410
rect 1170 680 1220 695
rect 1170 410 1185 680
rect 1205 410 1220 680
rect 1170 395 1220 410
rect 1270 680 1320 695
rect 1270 410 1285 680
rect 1305 410 1320 680
rect 1270 395 1320 410
<< ndiffc >>
rect 125 1780 145 2050
rect 225 1780 245 2050
rect 325 1780 345 2050
rect 425 1780 445 2050
rect 525 1780 545 2050
rect 625 1780 645 2050
rect 725 1780 745 2050
rect 825 1780 845 2050
rect 925 1780 945 2050
rect 1025 1780 1045 2050
rect 1125 1780 1145 2050
rect 125 1310 145 1580
rect 225 1310 245 1580
rect 325 1310 345 1580
rect 425 1310 445 1580
rect 525 1310 545 1580
rect 625 1310 645 1580
rect 725 1310 745 1580
rect 825 1310 845 1580
rect 925 1310 945 1580
rect 1025 1310 1045 1580
rect 1125 1310 1145 1580
rect -35 15 -15 285
rect 65 15 85 285
rect 165 15 185 285
rect 245 15 265 285
rect 345 15 365 285
rect 445 15 465 285
rect 525 15 545 285
rect 625 15 645 285
rect 725 15 745 285
rect 805 15 825 285
rect 905 15 925 285
rect 1005 15 1025 285
rect 1085 15 1105 285
rect 1185 15 1205 285
rect 1285 15 1305 285
rect 125 -390 145 -120
rect 225 -390 245 -120
rect 325 -390 345 -120
rect 425 -390 445 -120
rect 525 -390 545 -120
rect 625 -390 645 -120
rect 725 -390 745 -120
rect 825 -390 845 -120
rect 925 -390 945 -120
rect 1025 -390 1045 -120
rect 1125 -390 1145 -120
<< pdiffc >>
rect 125 830 145 1100
rect 225 830 245 1100
rect 325 830 345 1100
rect 425 830 445 1100
rect 525 830 545 1100
rect 625 830 645 1100
rect 725 830 745 1100
rect 825 830 845 1100
rect 925 830 945 1100
rect 1025 830 1045 1100
rect 1125 830 1145 1100
rect -35 410 -15 680
rect 65 410 85 680
rect 165 410 185 680
rect 245 410 265 680
rect 345 410 365 680
rect 445 410 465 680
rect 525 410 545 680
rect 625 410 645 680
rect 725 410 745 680
rect 805 410 825 680
rect 905 410 925 680
rect 1005 410 1025 680
rect 1085 410 1105 680
rect 1185 410 1205 680
rect 1285 410 1305 680
<< poly >>
rect 160 2110 210 2120
rect 160 2090 175 2110
rect 195 2090 210 2110
rect 160 2065 210 2090
rect 260 2080 1010 2130
rect 260 2065 310 2080
rect 360 2065 410 2080
rect 460 2065 510 2080
rect 560 2065 610 2080
rect 660 2065 710 2080
rect 760 2065 810 2080
rect 860 2065 910 2080
rect 960 2065 1010 2080
rect 1060 2110 1110 2120
rect 1060 2090 1075 2110
rect 1095 2090 1110 2110
rect 1060 2065 1110 2090
rect 160 1750 210 1765
rect 260 1750 310 1765
rect 360 1750 410 1765
rect 460 1750 510 1765
rect 560 1750 610 1765
rect 660 1750 710 1765
rect 760 1750 810 1765
rect 860 1750 910 1765
rect 960 1750 1010 1765
rect 1060 1750 1110 1765
rect 110 1685 285 1725
rect 110 1675 910 1685
rect 160 1640 210 1650
rect 160 1620 175 1640
rect 195 1620 210 1640
rect 235 1635 910 1675
rect 160 1595 210 1620
rect 260 1595 310 1610
rect 360 1595 410 1635
rect 460 1595 510 1635
rect 560 1595 610 1610
rect 660 1595 710 1610
rect 760 1595 810 1635
rect 860 1595 910 1635
rect 1060 1640 1110 1650
rect 1060 1620 1075 1640
rect 1095 1620 1110 1640
rect 960 1595 1010 1610
rect 1060 1595 1110 1620
rect 160 1280 210 1295
rect 260 1255 310 1295
rect 360 1280 410 1295
rect 460 1280 510 1295
rect 560 1255 610 1295
rect 660 1255 710 1295
rect 760 1280 810 1295
rect 860 1280 910 1295
rect 960 1255 1010 1295
rect 1060 1280 1110 1295
rect 110 1205 1010 1255
rect 160 1160 210 1170
rect 160 1140 175 1160
rect 195 1140 210 1160
rect 160 1115 210 1140
rect 260 1130 1010 1180
rect 260 1115 310 1130
rect 360 1115 410 1130
rect 460 1115 510 1130
rect 560 1115 610 1130
rect 660 1115 710 1130
rect 760 1115 810 1130
rect 860 1115 910 1130
rect 960 1115 1010 1130
rect 1060 1160 1110 1170
rect 1060 1140 1075 1160
rect 1095 1140 1110 1160
rect 1060 1115 1110 1140
rect 160 800 210 815
rect 260 800 310 815
rect 360 800 410 815
rect 460 800 510 815
rect 560 800 610 815
rect 660 800 710 815
rect 760 800 810 815
rect 860 800 910 815
rect 960 800 1010 815
rect 1060 800 1110 815
rect 0 740 50 750
rect 0 720 15 740
rect 35 720 50 740
rect 0 695 50 720
rect 100 710 1170 760
rect 100 695 150 710
rect 280 695 330 710
rect 380 695 430 710
rect 560 695 610 710
rect 660 695 710 710
rect 840 695 890 710
rect 940 695 990 710
rect 1120 695 1170 710
rect 1220 740 1270 750
rect 1220 720 1235 740
rect 1255 720 1270 740
rect 1220 695 1270 720
rect 0 380 50 395
rect 100 380 150 395
rect 280 380 330 395
rect 380 380 430 395
rect 560 380 610 395
rect 660 380 710 395
rect 840 380 890 395
rect 940 380 990 395
rect 1120 380 1170 395
rect 1220 380 1270 395
rect 475 345 805 355
rect 475 325 485 345
rect 505 340 775 345
rect 505 325 515 340
rect 475 315 515 325
rect 765 325 775 340
rect 795 325 805 345
rect 765 315 805 325
rect 0 300 50 315
rect 100 300 150 315
rect 280 300 330 315
rect 380 300 430 315
rect 560 300 610 315
rect 660 300 710 315
rect 840 300 890 315
rect 940 300 990 315
rect 1120 300 1170 315
rect 1220 300 1270 315
rect 0 -25 50 0
rect 0 -45 15 -25
rect 35 -45 50 -25
rect 0 -55 50 -45
rect 100 -15 150 0
rect 280 -15 330 0
rect 380 -15 430 0
rect 560 -15 610 0
rect 660 -15 710 0
rect 840 -15 890 0
rect 940 -15 990 0
rect 1120 -15 1170 0
rect 100 -65 1170 -15
rect 1220 -25 1270 0
rect 1220 -45 1235 -25
rect 1255 -45 1270 -25
rect 1220 -55 1270 -45
rect 160 -105 210 -90
rect 260 -105 310 -90
rect 360 -105 410 -90
rect 460 -105 510 -90
rect 560 -105 610 -90
rect 660 -105 710 -90
rect 760 -105 810 -90
rect 860 -105 910 -90
rect 960 -105 1010 -90
rect 1060 -105 1110 -90
rect 160 -430 210 -405
rect 160 -450 175 -430
rect 195 -450 210 -430
rect 160 -460 210 -450
rect 260 -420 310 -405
rect 360 -420 410 -405
rect 460 -420 510 -405
rect 560 -420 610 -405
rect 660 -420 710 -405
rect 760 -420 810 -405
rect 860 -420 910 -405
rect 960 -420 1010 -405
rect 260 -470 1010 -420
rect 1060 -430 1110 -405
rect 1060 -450 1075 -430
rect 1095 -450 1110 -430
rect 1060 -460 1110 -450
<< polycont >>
rect 175 2090 195 2110
rect 1075 2090 1095 2110
rect 175 1620 195 1640
rect 1075 1620 1095 1640
rect 175 1140 195 1160
rect 1075 1140 1095 1160
rect 15 720 35 740
rect 1235 720 1255 740
rect 485 325 505 345
rect 775 325 795 345
rect 15 -45 35 -25
rect 1235 -45 1255 -25
rect 175 -450 195 -430
rect 1075 -450 1095 -430
<< locali >>
rect 165 2110 205 2120
rect 165 2090 175 2110
rect 195 2090 205 2110
rect 165 2080 205 2090
rect 1065 2110 1105 2120
rect 1065 2090 1075 2110
rect 1095 2090 1105 2110
rect 1065 2080 1105 2090
rect 115 2050 155 2060
rect 115 1780 125 2050
rect 145 1780 155 2050
rect 115 1770 155 1780
rect 215 2050 255 2060
rect 215 1780 225 2050
rect 245 1780 255 2050
rect 215 1770 255 1780
rect 315 2050 355 2060
rect 315 1780 325 2050
rect 345 1780 355 2050
rect 315 1770 355 1780
rect 415 2050 455 2060
rect 415 1780 425 2050
rect 445 1780 455 2050
rect 415 1770 455 1780
rect 515 2050 555 2060
rect 515 1780 525 2050
rect 545 1780 555 2050
rect 515 1770 555 1780
rect 615 2050 655 2060
rect 615 1780 625 2050
rect 645 1780 655 2050
rect 615 1770 655 1780
rect 715 2050 755 2060
rect 715 1780 725 2050
rect 745 1780 755 2050
rect 715 1770 755 1780
rect 815 2050 855 2060
rect 815 1780 825 2050
rect 845 1780 855 2050
rect 815 1770 855 1780
rect 915 2050 955 2060
rect 915 1780 925 2050
rect 945 1780 955 2050
rect 915 1770 955 1780
rect 1015 2050 1055 2060
rect 1015 1780 1025 2050
rect 1045 1780 1055 2050
rect 1015 1770 1055 1780
rect 1115 2050 1155 2060
rect 1115 1780 1125 2050
rect 1145 1780 1155 2050
rect 1115 1770 1155 1780
rect 235 1690 255 1770
rect 425 1690 445 1770
rect 625 1690 645 1770
rect 825 1690 845 1770
rect 1015 1690 1035 1770
rect 235 1670 1035 1690
rect 165 1640 205 1650
rect 165 1620 175 1640
rect 195 1620 205 1640
rect 165 1610 205 1620
rect 325 1590 345 1670
rect 525 1590 545 1670
rect 725 1590 745 1670
rect 925 1590 945 1670
rect 1065 1640 1105 1650
rect 1065 1620 1075 1640
rect 1095 1620 1105 1640
rect 1065 1610 1105 1620
rect 115 1580 155 1590
rect 115 1310 125 1580
rect 145 1310 155 1580
rect 115 1300 155 1310
rect 215 1580 255 1590
rect 215 1310 225 1580
rect 245 1310 255 1580
rect 215 1300 255 1310
rect 315 1580 355 1590
rect 315 1310 325 1580
rect 345 1310 355 1580
rect 315 1300 355 1310
rect 415 1580 455 1590
rect 415 1310 425 1580
rect 445 1310 455 1580
rect 415 1300 455 1310
rect 515 1580 555 1590
rect 515 1310 525 1580
rect 545 1310 555 1580
rect 515 1300 555 1310
rect 615 1580 655 1590
rect 615 1310 625 1580
rect 645 1310 655 1580
rect 615 1300 655 1310
rect 715 1580 755 1590
rect 715 1310 725 1580
rect 745 1310 755 1580
rect 715 1300 755 1310
rect 815 1580 855 1590
rect 815 1310 825 1580
rect 845 1310 855 1580
rect 815 1300 855 1310
rect 915 1580 955 1590
rect 915 1310 925 1580
rect 945 1310 955 1580
rect 915 1300 955 1310
rect 1015 1580 1055 1590
rect 1015 1310 1025 1580
rect 1045 1310 1055 1580
rect 1015 1300 1055 1310
rect 1115 1580 1155 1590
rect 1115 1310 1125 1580
rect 1145 1310 1155 1580
rect 1115 1300 1155 1310
rect 165 1160 205 1170
rect 165 1140 175 1160
rect 195 1140 205 1160
rect 165 1130 205 1140
rect 225 1110 245 1300
rect 425 1110 445 1300
rect 625 1110 645 1300
rect 825 1110 845 1300
rect 1025 1110 1045 1300
rect 1065 1160 1105 1170
rect 1065 1140 1075 1160
rect 1095 1140 1105 1160
rect 1065 1130 1105 1140
rect 115 1100 155 1110
rect 115 830 125 1100
rect 145 830 155 1100
rect 115 820 155 830
rect 215 1100 255 1110
rect 215 830 225 1100
rect 245 830 255 1100
rect 215 820 255 830
rect 315 1100 355 1110
rect 315 830 325 1100
rect 345 830 355 1100
rect 315 820 355 830
rect 415 1100 455 1110
rect 415 830 425 1100
rect 445 830 455 1100
rect 415 820 455 830
rect 515 1100 555 1110
rect 515 830 525 1100
rect 545 830 555 1100
rect 515 820 555 830
rect 615 1100 655 1110
rect 615 830 625 1100
rect 645 830 655 1100
rect 615 820 655 830
rect 715 1100 755 1110
rect 715 830 725 1100
rect 745 830 755 1100
rect 715 820 755 830
rect 815 1100 855 1110
rect 815 830 825 1100
rect 845 830 855 1100
rect 815 820 855 830
rect 915 1100 955 1110
rect 915 830 925 1100
rect 945 830 955 1100
rect 915 820 955 830
rect 1015 1100 1055 1110
rect 1015 830 1025 1100
rect 1045 830 1055 1100
rect 1015 820 1055 830
rect 1115 1100 1155 1110
rect 1115 830 1125 1100
rect 1145 830 1155 1100
rect 1115 820 1155 830
rect 225 800 245 820
rect 425 800 445 820
rect 625 800 645 820
rect 825 800 845 820
rect 1025 800 1045 820
rect 5 740 45 750
rect 5 720 15 740
rect 35 720 45 740
rect 5 710 45 720
rect 1225 740 1265 750
rect 1225 720 1235 740
rect 1255 720 1265 740
rect 1225 710 1265 720
rect 65 690 85 710
rect 345 690 365 700
rect 625 690 645 700
rect 905 690 925 700
rect 1185 690 1205 700
rect -45 680 -5 690
rect -45 410 -35 680
rect -15 410 -5 680
rect -45 400 -5 410
rect 55 680 95 690
rect 55 410 65 680
rect 85 410 95 680
rect 55 400 95 410
rect 155 680 195 690
rect 155 410 165 680
rect 185 410 195 680
rect 155 400 195 410
rect 235 680 275 690
rect 235 410 245 680
rect 265 410 275 680
rect 235 400 275 410
rect 335 680 375 690
rect 335 410 345 680
rect 365 410 375 680
rect 335 400 375 410
rect 435 680 475 690
rect 435 410 445 680
rect 465 410 475 680
rect 435 400 475 410
rect 515 680 555 690
rect 515 410 525 680
rect 545 410 555 680
rect 515 400 555 410
rect 615 680 655 690
rect 615 410 625 680
rect 645 410 655 680
rect 615 400 655 410
rect 715 680 755 690
rect 715 410 725 680
rect 745 410 755 680
rect 715 400 755 410
rect 795 680 835 690
rect 795 410 805 680
rect 825 410 835 680
rect 795 400 835 410
rect 895 680 935 690
rect 895 410 905 680
rect 925 410 935 680
rect 895 400 935 410
rect 995 680 1035 690
rect 995 410 1005 680
rect 1025 410 1035 680
rect 995 400 1035 410
rect 1075 680 1115 690
rect 1075 410 1085 680
rect 1105 410 1115 680
rect 1075 400 1115 410
rect 1175 680 1215 690
rect 1175 410 1185 680
rect 1205 410 1215 680
rect 1175 400 1215 410
rect 1275 680 1315 690
rect 1275 410 1285 680
rect 1305 410 1315 680
rect 1275 400 1315 410
rect 175 355 195 400
rect 175 345 215 355
rect 175 325 185 345
rect 205 325 215 345
rect 175 315 215 325
rect 245 335 265 400
rect 455 355 475 400
rect 455 345 515 355
rect 455 335 485 345
rect 245 325 485 335
rect 505 325 515 345
rect 245 315 515 325
rect 535 335 555 400
rect 615 345 655 355
rect 615 335 625 345
rect 535 325 625 335
rect 645 335 655 345
rect 725 335 745 400
rect 805 355 825 400
rect 645 325 745 335
rect 535 315 745 325
rect 765 345 825 355
rect 765 325 775 345
rect 795 335 825 345
rect 1005 335 1025 400
rect 1075 355 1095 400
rect 795 325 1025 335
rect 765 315 1025 325
rect 1055 345 1095 355
rect 1055 325 1065 345
rect 1085 325 1095 345
rect 1055 315 1095 325
rect 175 295 195 315
rect 245 295 265 315
rect 455 295 475 315
rect 535 295 555 315
rect 725 295 745 315
rect 805 295 825 315
rect 1005 295 1025 315
rect 1075 295 1095 315
rect -45 285 -5 295
rect -45 15 -35 285
rect -15 15 -5 285
rect -45 5 -5 15
rect 55 285 95 295
rect 55 15 65 285
rect 85 15 95 285
rect 55 5 95 15
rect 155 285 195 295
rect 155 15 165 285
rect 185 15 195 285
rect 155 5 195 15
rect 235 285 275 295
rect 235 15 245 285
rect 265 15 275 285
rect 235 5 275 15
rect 335 285 375 295
rect 335 15 345 285
rect 365 15 375 285
rect 335 5 375 15
rect 435 285 475 295
rect 435 15 445 285
rect 465 15 475 285
rect 435 5 475 15
rect 515 285 555 295
rect 515 15 525 285
rect 545 15 555 285
rect 515 5 555 15
rect 615 285 655 295
rect 615 15 625 285
rect 645 15 655 285
rect 615 5 655 15
rect 715 285 755 295
rect 715 15 725 285
rect 745 15 755 285
rect 715 5 755 15
rect 795 285 835 295
rect 795 15 805 285
rect 825 15 835 285
rect 795 5 835 15
rect 895 285 935 295
rect 895 15 905 285
rect 925 15 935 285
rect 895 5 935 15
rect 995 285 1035 295
rect 995 15 1005 285
rect 1025 15 1035 285
rect 995 5 1035 15
rect 1075 285 1115 295
rect 1075 15 1085 285
rect 1105 15 1115 285
rect 1075 5 1115 15
rect 1175 285 1215 295
rect 1175 15 1185 285
rect 1205 15 1215 285
rect 1175 5 1215 15
rect 1275 285 1315 295
rect 1275 15 1285 285
rect 1305 15 1315 285
rect 1275 5 1315 15
rect 5 -25 45 -15
rect 5 -45 15 -25
rect 35 -45 45 -25
rect 5 -55 45 -45
rect 65 -70 85 5
rect 345 -70 365 5
rect 225 -110 245 -75
rect 425 -110 445 -70
rect 625 -110 645 5
rect 905 -75 925 5
rect 1185 -75 1205 5
rect 1225 -25 1265 -15
rect 1225 -45 1235 -25
rect 1255 -45 1265 -25
rect 1225 -55 1265 -45
rect 825 -110 845 -75
rect 1025 -110 1045 -75
rect 115 -120 155 -110
rect 115 -390 125 -120
rect 145 -390 155 -120
rect 115 -400 155 -390
rect 215 -120 255 -110
rect 215 -390 225 -120
rect 245 -390 255 -120
rect 215 -400 255 -390
rect 315 -120 355 -110
rect 315 -390 325 -120
rect 345 -390 355 -120
rect 315 -400 355 -390
rect 415 -120 455 -110
rect 415 -390 425 -120
rect 445 -390 455 -120
rect 415 -400 455 -390
rect 515 -120 555 -110
rect 515 -390 525 -120
rect 545 -390 555 -120
rect 515 -400 555 -390
rect 615 -120 655 -110
rect 615 -390 625 -120
rect 645 -390 655 -120
rect 615 -400 655 -390
rect 715 -120 755 -110
rect 715 -390 725 -120
rect 745 -390 755 -120
rect 715 -400 755 -390
rect 815 -120 855 -110
rect 815 -390 825 -120
rect 845 -390 855 -120
rect 815 -400 855 -390
rect 915 -120 955 -110
rect 915 -390 925 -120
rect 945 -390 955 -120
rect 915 -400 955 -390
rect 1015 -120 1055 -110
rect 1015 -390 1025 -120
rect 1045 -390 1055 -120
rect 1015 -400 1055 -390
rect 1115 -120 1155 -110
rect 1115 -390 1125 -120
rect 1145 -390 1155 -120
rect 1115 -400 1155 -390
rect 165 -430 205 -420
rect 165 -450 175 -430
rect 195 -450 205 -430
rect 165 -460 205 -450
rect 1065 -430 1105 -420
rect 1065 -450 1075 -430
rect 1095 -450 1105 -430
rect 1065 -460 1105 -450
<< viali >>
rect 125 1780 145 2050
rect 325 1780 345 2050
rect 525 1780 545 2050
rect 725 1780 745 2050
rect 925 1780 945 2050
rect 1125 1780 1145 2050
rect 125 1310 145 1580
rect 1125 1310 1145 1580
rect 125 830 145 1100
rect 325 830 345 1100
rect 525 830 545 1100
rect 725 830 745 1100
rect 925 830 945 1100
rect 1125 830 1145 1100
rect 185 325 205 345
rect 625 325 645 345
rect 1065 325 1085 345
rect 125 -390 145 -120
rect 325 -390 345 -120
rect 525 -390 545 -120
rect 725 -390 745 -120
rect 925 -390 945 -120
rect 1125 -390 1145 -120
<< metal1 >>
rect 175 345 1095 355
rect 175 325 185 345
rect 205 340 625 345
rect 205 325 215 340
rect 175 315 215 325
rect 615 325 625 340
rect 645 340 1065 345
rect 645 325 655 340
rect 615 315 655 325
rect 1055 325 1065 340
rect 1085 325 1095 345
rect 1055 315 1095 325
<< end >>
