magic
tech sky130A
timestamp 1697083663
<< error_p >>
rect 125 2062 145 2065
rect 125 1798 128 2062
rect 142 1798 145 2062
rect 125 1795 145 1798
rect 325 2062 345 2065
rect 325 1798 328 2062
rect 342 1798 345 2062
rect 325 1795 345 1798
rect 525 2062 545 2065
rect 525 1798 528 2062
rect 542 1798 545 2062
rect 525 1795 545 1798
rect 725 2062 745 2065
rect 725 1798 728 2062
rect 742 1798 745 2062
rect 725 1795 745 1798
rect 925 2062 945 2065
rect 925 1798 928 2062
rect 942 1798 945 2062
rect 925 1795 945 1798
rect 1125 2062 1145 2065
rect 1125 1798 1128 2062
rect 1142 1798 1145 2062
rect 1125 1795 1145 1798
rect 125 1627 145 1630
rect 125 1363 128 1627
rect 142 1363 145 1627
rect 125 1360 145 1363
rect 1125 1627 1145 1630
rect 1125 1363 1128 1627
rect 1142 1363 1145 1627
rect 1125 1360 1145 1363
rect 125 1122 145 1125
rect 125 858 128 1122
rect 142 858 145 1122
rect 125 855 145 858
rect 325 1122 345 1125
rect 325 858 328 1122
rect 342 858 345 1122
rect 325 855 345 858
rect 525 1122 545 1125
rect 525 858 528 1122
rect 542 858 545 1122
rect 525 855 545 858
rect 725 1122 745 1125
rect 725 858 728 1122
rect 742 858 745 1122
rect 725 855 745 858
rect 925 1122 945 1125
rect 925 858 928 1122
rect 942 858 945 1122
rect 925 855 945 858
rect 1125 1122 1145 1125
rect 1125 858 1128 1122
rect 1142 858 1145 1122
rect 1125 855 1145 858
rect 125 -83 145 -80
rect 125 -347 128 -83
rect 142 -347 145 -83
rect 125 -350 145 -347
rect 325 -83 345 -80
rect 325 -347 328 -83
rect 342 -347 345 -83
rect 325 -350 345 -347
rect 525 -83 545 -80
rect 525 -347 528 -83
rect 542 -347 545 -83
rect 525 -350 545 -347
rect 725 -83 745 -80
rect 725 -347 728 -83
rect 742 -347 745 -83
rect 725 -350 745 -347
rect 925 -83 945 -80
rect 925 -347 928 -83
rect 942 -347 945 -83
rect 925 -350 945 -347
rect 1125 -83 1145 -80
rect 1125 -347 1128 -83
rect 1142 -347 1145 -83
rect 1125 -350 1145 -347
<< nwell >>
rect 90 775 1180 1160
rect -70 375 1340 775
<< nmos >>
rect 160 1780 210 2080
rect 260 1780 310 2080
rect 360 1780 410 2080
rect 460 1780 510 2080
rect 560 1780 610 2080
rect 660 1780 710 2080
rect 760 1780 810 2080
rect 860 1780 910 2080
rect 960 1780 1010 2080
rect 1060 1780 1110 2080
rect 160 1345 210 1645
rect 260 1345 310 1645
rect 360 1345 410 1645
rect 460 1345 510 1645
rect 560 1345 610 1645
rect 660 1345 710 1645
rect 760 1345 810 1645
rect 860 1345 910 1645
rect 960 1345 1010 1645
rect 1060 1345 1110 1645
rect 0 40 50 340
rect 100 40 150 340
rect 280 40 330 340
rect 380 40 430 340
rect 560 40 610 340
rect 660 40 710 340
rect 840 40 890 340
rect 940 40 990 340
rect 1120 40 1170 340
rect 1220 40 1270 340
rect 160 -365 210 -65
rect 260 -365 310 -65
rect 360 -365 410 -65
rect 460 -365 510 -65
rect 560 -365 610 -65
rect 660 -365 710 -65
rect 760 -365 810 -65
rect 860 -365 910 -65
rect 960 -365 1010 -65
rect 1060 -365 1110 -65
<< pmos >>
rect 160 840 210 1140
rect 260 840 310 1140
rect 360 840 410 1140
rect 460 840 510 1140
rect 560 840 610 1140
rect 660 840 710 1140
rect 760 840 810 1140
rect 860 840 910 1140
rect 960 840 1010 1140
rect 1060 840 1110 1140
rect 0 395 50 695
rect 100 395 150 695
rect 280 395 330 695
rect 380 395 430 695
rect 560 395 610 695
rect 660 395 710 695
rect 840 395 890 695
rect 940 395 990 695
rect 1120 395 1170 695
rect 1220 395 1270 695
<< ndiff >>
rect 110 2065 160 2080
rect 110 1795 125 2065
rect 145 1795 160 2065
rect 110 1780 160 1795
rect 210 2065 260 2080
rect 210 1795 225 2065
rect 245 1795 260 2065
rect 210 1780 260 1795
rect 310 2065 360 2080
rect 310 1795 325 2065
rect 345 1795 360 2065
rect 310 1780 360 1795
rect 410 2065 460 2080
rect 410 1795 425 2065
rect 445 1795 460 2065
rect 410 1780 460 1795
rect 510 2065 560 2080
rect 510 1795 525 2065
rect 545 1795 560 2065
rect 510 1780 560 1795
rect 610 2065 660 2080
rect 610 1795 625 2065
rect 645 1795 660 2065
rect 610 1780 660 1795
rect 710 2065 760 2080
rect 710 1795 725 2065
rect 745 1795 760 2065
rect 710 1780 760 1795
rect 810 2065 860 2080
rect 810 1795 825 2065
rect 845 1795 860 2065
rect 810 1780 860 1795
rect 910 2065 960 2080
rect 910 1795 925 2065
rect 945 1795 960 2065
rect 910 1780 960 1795
rect 1010 2065 1060 2080
rect 1010 1795 1025 2065
rect 1045 1795 1060 2065
rect 1010 1780 1060 1795
rect 1110 2065 1160 2080
rect 1110 1795 1125 2065
rect 1145 1795 1160 2065
rect 1110 1780 1160 1795
rect 110 1630 160 1645
rect 110 1360 125 1630
rect 145 1360 160 1630
rect 110 1345 160 1360
rect 210 1630 260 1645
rect 210 1360 225 1630
rect 245 1360 260 1630
rect 210 1345 260 1360
rect 310 1630 360 1645
rect 310 1360 325 1630
rect 345 1360 360 1630
rect 310 1345 360 1360
rect 410 1630 460 1645
rect 410 1360 425 1630
rect 445 1360 460 1630
rect 410 1345 460 1360
rect 510 1630 560 1645
rect 510 1360 525 1630
rect 545 1360 560 1630
rect 510 1345 560 1360
rect 610 1630 660 1645
rect 610 1360 625 1630
rect 645 1360 660 1630
rect 610 1345 660 1360
rect 710 1630 760 1645
rect 710 1360 725 1630
rect 745 1360 760 1630
rect 710 1345 760 1360
rect 810 1630 860 1645
rect 810 1360 825 1630
rect 845 1360 860 1630
rect 810 1345 860 1360
rect 910 1630 960 1645
rect 910 1360 925 1630
rect 945 1360 960 1630
rect 910 1345 960 1360
rect 1010 1630 1060 1645
rect 1010 1360 1025 1630
rect 1045 1360 1060 1630
rect 1010 1345 1060 1360
rect 1110 1630 1160 1645
rect 1110 1360 1125 1630
rect 1145 1360 1160 1630
rect 1110 1345 1160 1360
rect -50 325 0 340
rect -50 55 -35 325
rect -15 55 0 325
rect -50 40 0 55
rect 50 325 100 340
rect 50 55 65 325
rect 85 55 100 325
rect 50 40 100 55
rect 150 325 200 340
rect 150 55 165 325
rect 185 55 200 325
rect 150 40 200 55
rect 230 325 280 340
rect 230 55 245 325
rect 265 55 280 325
rect 230 40 280 55
rect 330 325 380 340
rect 330 55 345 325
rect 365 55 380 325
rect 330 40 380 55
rect 430 325 480 340
rect 430 55 445 325
rect 465 55 480 325
rect 430 40 480 55
rect 510 325 560 340
rect 510 55 525 325
rect 545 55 560 325
rect 510 40 560 55
rect 610 325 660 340
rect 610 55 625 325
rect 645 55 660 325
rect 610 40 660 55
rect 710 325 760 340
rect 710 55 725 325
rect 745 55 760 325
rect 710 40 760 55
rect 790 325 840 340
rect 790 55 805 325
rect 825 55 840 325
rect 790 40 840 55
rect 890 325 940 340
rect 890 55 905 325
rect 925 55 940 325
rect 890 40 940 55
rect 990 325 1040 340
rect 990 55 1005 325
rect 1025 55 1040 325
rect 990 40 1040 55
rect 1070 325 1120 340
rect 1070 55 1085 325
rect 1105 55 1120 325
rect 1070 40 1120 55
rect 1170 325 1220 340
rect 1170 55 1185 325
rect 1205 55 1220 325
rect 1170 40 1220 55
rect 1270 325 1320 340
rect 1270 55 1285 325
rect 1305 55 1320 325
rect 1270 40 1320 55
rect 110 -80 160 -65
rect 110 -350 125 -80
rect 145 -350 160 -80
rect 110 -365 160 -350
rect 210 -80 260 -65
rect 210 -350 225 -80
rect 245 -350 260 -80
rect 210 -365 260 -350
rect 310 -80 360 -65
rect 310 -350 325 -80
rect 345 -350 360 -80
rect 310 -365 360 -350
rect 410 -80 460 -65
rect 410 -350 425 -80
rect 445 -350 460 -80
rect 410 -365 460 -350
rect 510 -80 560 -65
rect 510 -350 525 -80
rect 545 -350 560 -80
rect 510 -365 560 -350
rect 610 -80 660 -65
rect 610 -350 625 -80
rect 645 -350 660 -80
rect 610 -365 660 -350
rect 710 -80 760 -65
rect 710 -350 725 -80
rect 745 -350 760 -80
rect 710 -365 760 -350
rect 810 -80 860 -65
rect 810 -350 825 -80
rect 845 -350 860 -80
rect 810 -365 860 -350
rect 910 -80 960 -65
rect 910 -350 925 -80
rect 945 -350 960 -80
rect 910 -365 960 -350
rect 1010 -80 1060 -65
rect 1010 -350 1025 -80
rect 1045 -350 1060 -80
rect 1010 -365 1060 -350
rect 1110 -80 1160 -65
rect 1110 -350 1125 -80
rect 1145 -350 1160 -80
rect 1110 -365 1160 -350
<< pdiff >>
rect 110 1125 160 1140
rect 110 855 125 1125
rect 145 855 160 1125
rect 110 840 160 855
rect 210 1125 260 1140
rect 210 855 225 1125
rect 245 855 260 1125
rect 210 840 260 855
rect 310 1125 360 1140
rect 310 855 325 1125
rect 345 855 360 1125
rect 310 840 360 855
rect 410 1125 460 1140
rect 410 855 425 1125
rect 445 855 460 1125
rect 410 840 460 855
rect 510 1125 560 1140
rect 510 855 525 1125
rect 545 855 560 1125
rect 510 840 560 855
rect 610 1125 660 1140
rect 610 855 625 1125
rect 645 855 660 1125
rect 610 840 660 855
rect 710 1125 760 1140
rect 710 855 725 1125
rect 745 855 760 1125
rect 710 840 760 855
rect 810 1125 860 1140
rect 810 855 825 1125
rect 845 855 860 1125
rect 810 840 860 855
rect 910 1125 960 1140
rect 910 855 925 1125
rect 945 855 960 1125
rect 910 840 960 855
rect 1010 1125 1060 1140
rect 1010 855 1025 1125
rect 1045 855 1060 1125
rect 1010 840 1060 855
rect 1110 1125 1160 1140
rect 1110 855 1125 1125
rect 1145 855 1160 1125
rect 1110 840 1160 855
rect -50 680 0 695
rect -50 410 -35 680
rect -15 410 0 680
rect -50 395 0 410
rect 50 680 100 695
rect 50 410 65 680
rect 85 410 100 680
rect 50 395 100 410
rect 150 680 200 695
rect 150 410 165 680
rect 185 410 200 680
rect 150 395 200 410
rect 230 680 280 695
rect 230 410 245 680
rect 265 410 280 680
rect 230 395 280 410
rect 330 680 380 695
rect 330 410 345 680
rect 365 410 380 680
rect 330 395 380 410
rect 430 680 480 695
rect 430 410 445 680
rect 465 410 480 680
rect 430 395 480 410
rect 510 680 560 695
rect 510 410 525 680
rect 545 410 560 680
rect 510 395 560 410
rect 610 680 660 695
rect 610 410 625 680
rect 645 410 660 680
rect 610 395 660 410
rect 710 680 760 695
rect 710 410 725 680
rect 745 410 760 680
rect 710 395 760 410
rect 790 680 840 695
rect 790 410 805 680
rect 825 410 840 680
rect 790 395 840 410
rect 890 680 940 695
rect 890 410 905 680
rect 925 410 940 680
rect 890 395 940 410
rect 990 680 1040 695
rect 990 410 1005 680
rect 1025 410 1040 680
rect 990 395 1040 410
rect 1070 680 1120 695
rect 1070 410 1085 680
rect 1105 410 1120 680
rect 1070 395 1120 410
rect 1170 680 1220 695
rect 1170 410 1185 680
rect 1205 410 1220 680
rect 1170 395 1220 410
rect 1270 680 1320 695
rect 1270 410 1285 680
rect 1305 410 1320 680
rect 1270 395 1320 410
<< ndiffc >>
rect 125 1795 145 2065
rect 225 1795 245 2065
rect 325 1795 345 2065
rect 425 1795 445 2065
rect 525 1795 545 2065
rect 625 1795 645 2065
rect 725 1795 745 2065
rect 825 1795 845 2065
rect 925 1795 945 2065
rect 1025 1795 1045 2065
rect 1125 1795 1145 2065
rect 125 1360 145 1630
rect 225 1360 245 1630
rect 325 1360 345 1630
rect 425 1360 445 1630
rect 525 1360 545 1630
rect 625 1360 645 1630
rect 725 1360 745 1630
rect 825 1360 845 1630
rect 925 1360 945 1630
rect 1025 1360 1045 1630
rect 1125 1360 1145 1630
rect -35 55 -15 325
rect 65 55 85 325
rect 165 55 185 325
rect 245 55 265 325
rect 345 55 365 325
rect 445 55 465 325
rect 525 55 545 325
rect 625 55 645 325
rect 725 55 745 325
rect 805 55 825 325
rect 905 55 925 325
rect 1005 55 1025 325
rect 1085 55 1105 325
rect 1185 55 1205 325
rect 1285 55 1305 325
rect 125 -350 145 -80
rect 225 -350 245 -80
rect 325 -350 345 -80
rect 425 -350 445 -80
rect 525 -350 545 -80
rect 625 -350 645 -80
rect 725 -350 745 -80
rect 825 -350 845 -80
rect 925 -350 945 -80
rect 1025 -350 1045 -80
rect 1125 -350 1145 -80
<< pdiffc >>
rect 125 855 145 1125
rect 225 855 245 1125
rect 325 855 345 1125
rect 425 855 445 1125
rect 525 855 545 1125
rect 625 855 645 1125
rect 725 855 745 1125
rect 825 855 845 1125
rect 925 855 945 1125
rect 1025 855 1045 1125
rect 1125 855 1145 1125
rect -35 410 -15 680
rect 65 410 85 680
rect 165 410 185 680
rect 245 410 265 680
rect 345 410 365 680
rect 445 410 465 680
rect 525 410 545 680
rect 625 410 645 680
rect 725 410 745 680
rect 805 410 825 680
rect 905 410 925 680
rect 1005 410 1025 680
rect 1085 410 1105 680
rect 1185 410 1205 680
rect 1285 410 1305 680
<< poly >>
rect 160 2125 210 2135
rect 160 2105 175 2125
rect 195 2105 210 2125
rect 160 2080 210 2105
rect 260 2125 1010 2145
rect 260 2105 275 2125
rect 295 2105 1010 2125
rect 260 2095 1010 2105
rect 260 2080 310 2095
rect 360 2080 410 2095
rect 460 2080 510 2095
rect 560 2080 610 2095
rect 660 2080 710 2095
rect 760 2080 810 2095
rect 860 2080 910 2095
rect 960 2080 1010 2095
rect 1060 2125 1110 2135
rect 1060 2105 1075 2125
rect 1095 2105 1110 2125
rect 1060 2080 1110 2105
rect 160 1765 210 1780
rect 260 1765 310 1780
rect 360 1765 410 1780
rect 460 1765 510 1780
rect 560 1765 610 1780
rect 660 1765 710 1780
rect 760 1765 810 1780
rect 860 1765 910 1780
rect 960 1765 1010 1780
rect 1060 1765 1110 1780
rect 235 1715 910 1735
rect 160 1690 210 1700
rect 160 1670 175 1690
rect 195 1670 210 1690
rect 235 1695 245 1715
rect 265 1695 910 1715
rect 235 1685 910 1695
rect 160 1645 210 1670
rect 260 1645 310 1660
rect 360 1645 410 1685
rect 460 1645 510 1685
rect 560 1645 610 1660
rect 660 1645 710 1660
rect 760 1645 810 1685
rect 860 1645 910 1685
rect 1060 1690 1110 1700
rect 1060 1670 1075 1690
rect 1095 1670 1110 1690
rect 960 1645 1010 1660
rect 1060 1645 1110 1670
rect 160 1330 210 1345
rect 260 1305 310 1345
rect 360 1330 410 1345
rect 460 1330 510 1345
rect 560 1305 610 1345
rect 660 1305 710 1345
rect 760 1330 810 1345
rect 860 1330 910 1345
rect 960 1305 1010 1345
rect 1060 1330 1110 1345
rect 110 1255 1010 1305
rect 110 1205 310 1230
rect 110 1180 1010 1205
rect 260 1155 1010 1180
rect 160 1140 210 1155
rect 260 1140 310 1155
rect 360 1140 410 1155
rect 460 1140 510 1155
rect 560 1140 610 1155
rect 660 1140 710 1155
rect 760 1140 810 1155
rect 860 1140 910 1155
rect 960 1140 1010 1155
rect 1060 1140 1110 1155
rect -55 775 125 825
rect 160 815 210 840
rect 260 825 310 840
rect 360 825 410 840
rect 460 825 510 840
rect 560 825 610 840
rect 660 825 710 840
rect 760 825 810 840
rect 860 825 910 840
rect 960 825 1010 840
rect 160 795 175 815
rect 195 795 210 815
rect 160 785 210 795
rect 1060 815 1110 840
rect 1060 795 1075 815
rect 1095 795 1110 815
rect 1060 785 1110 795
rect 75 760 125 775
rect 0 740 50 750
rect 0 720 15 740
rect 35 720 50 740
rect 0 695 50 720
rect 75 710 1170 760
rect 100 695 150 710
rect 280 695 330 710
rect 380 695 430 710
rect 560 695 610 710
rect 660 695 710 710
rect 840 695 890 710
rect 940 695 990 710
rect 1120 695 1170 710
rect 1220 740 1270 750
rect 1220 720 1235 740
rect 1255 720 1270 740
rect 1220 695 1270 720
rect 0 380 50 395
rect 100 380 150 395
rect 280 380 330 395
rect 380 380 430 395
rect 560 380 610 395
rect 660 380 710 395
rect 840 380 890 395
rect 940 380 990 395
rect 1120 380 1170 395
rect 1220 380 1270 395
rect 0 340 50 355
rect 100 340 150 355
rect 280 340 330 355
rect 380 340 430 355
rect 560 340 610 355
rect 660 340 710 355
rect 840 340 890 355
rect 940 340 990 355
rect 1120 340 1170 355
rect 1220 340 1270 355
rect 0 15 50 40
rect 0 -5 15 15
rect 35 -5 50 15
rect 0 -15 50 -5
rect 100 25 150 40
rect 280 25 330 40
rect 380 25 430 40
rect 560 25 610 40
rect 660 25 710 40
rect 840 25 890 40
rect 940 25 990 40
rect 1120 25 1170 40
rect 100 15 1170 25
rect 100 -5 115 15
rect 135 -5 1170 15
rect 100 -25 1170 -5
rect 1220 15 1270 40
rect 1220 -5 1235 15
rect 1255 -5 1270 15
rect 1220 -15 1270 -5
rect 160 -65 210 -50
rect 260 -65 310 -50
rect 360 -65 410 -50
rect 460 -65 510 -50
rect 560 -65 610 -50
rect 660 -65 710 -50
rect 760 -65 810 -50
rect 860 -65 910 -50
rect 960 -65 1010 -50
rect 1060 -65 1110 -50
rect 160 -390 210 -365
rect 160 -410 175 -390
rect 195 -410 210 -390
rect 160 -420 210 -410
rect 260 -380 310 -365
rect 360 -380 410 -365
rect 460 -380 510 -365
rect 560 -380 610 -365
rect 660 -380 710 -365
rect 760 -380 810 -365
rect 860 -380 910 -365
rect 960 -380 1010 -365
rect 260 -430 1010 -380
rect 1060 -390 1110 -365
rect 1060 -410 1075 -390
rect 1095 -410 1110 -390
rect 1060 -420 1110 -410
<< polycont >>
rect 175 2105 195 2125
rect 275 2105 295 2125
rect 1075 2105 1095 2125
rect 175 1670 195 1690
rect 245 1695 265 1715
rect 1075 1670 1095 1690
rect 175 795 195 815
rect 1075 795 1095 815
rect 15 720 35 740
rect 1235 720 1255 740
rect 15 -5 35 15
rect 115 -5 135 15
rect 1235 -5 1255 15
rect 175 -410 195 -390
rect 1075 -410 1095 -390
<< locali >>
rect 120 2155 285 2175
rect 265 2135 285 2155
rect 165 2125 205 2135
rect 165 2105 175 2125
rect 195 2105 205 2125
rect 165 2095 205 2105
rect 265 2125 305 2135
rect 265 2105 275 2125
rect 295 2105 305 2125
rect 265 2095 305 2105
rect 1065 2125 1105 2135
rect 1065 2105 1075 2125
rect 1095 2105 1105 2125
rect 1065 2095 1105 2105
rect 115 2065 155 2075
rect 115 1795 125 2065
rect 145 1795 155 2065
rect 115 1785 155 1795
rect 215 2065 255 2075
rect 215 1795 225 2065
rect 245 1805 255 2065
rect 315 2065 355 2075
rect 245 1795 295 1805
rect 215 1785 295 1795
rect 315 1795 325 2065
rect 345 1795 355 2065
rect 315 1785 355 1795
rect 415 2065 455 2075
rect 415 1795 425 2065
rect 445 1795 455 2065
rect 415 1785 455 1795
rect 515 2065 555 2075
rect 515 1795 525 2065
rect 545 1795 555 2065
rect 515 1785 555 1795
rect 615 2065 655 2075
rect 615 1795 625 2065
rect 645 1795 655 2065
rect 615 1785 655 1795
rect 715 2065 755 2075
rect 715 1795 725 2065
rect 745 1795 755 2065
rect 715 1785 755 1795
rect 815 2065 855 2075
rect 815 1795 825 2065
rect 845 1795 855 2065
rect 815 1785 855 1795
rect 915 2065 955 2075
rect 915 1795 925 2065
rect 945 1795 955 2065
rect 915 1785 955 1795
rect 1015 2065 1055 2075
rect 1015 1795 1025 2065
rect 1045 1795 1055 2065
rect 1015 1785 1055 1795
rect 1115 2065 1155 2075
rect 1115 1795 1125 2065
rect 1145 1795 1155 2065
rect 1115 1785 1155 1795
rect 275 1765 295 1785
rect 275 1745 345 1765
rect 110 1725 255 1745
rect 325 1740 345 1745
rect 425 1740 445 1785
rect 625 1740 645 1785
rect 825 1740 845 1785
rect 1015 1740 1035 1785
rect 235 1715 275 1725
rect 165 1690 205 1700
rect 165 1670 175 1690
rect 195 1670 205 1690
rect 235 1695 245 1715
rect 265 1695 275 1715
rect 235 1685 275 1695
rect 325 1720 1035 1740
rect 165 1660 205 1670
rect 325 1640 345 1720
rect 525 1640 545 1720
rect 725 1640 745 1720
rect 925 1640 945 1720
rect 1065 1690 1105 1700
rect 1065 1670 1075 1690
rect 1095 1670 1105 1690
rect 1065 1660 1105 1670
rect 115 1630 155 1640
rect 115 1360 125 1630
rect 145 1360 155 1630
rect 115 1350 155 1360
rect 215 1630 255 1640
rect 215 1360 225 1630
rect 245 1360 255 1630
rect 215 1350 255 1360
rect 315 1630 355 1640
rect 315 1360 325 1630
rect 345 1360 355 1630
rect 315 1350 355 1360
rect 415 1630 455 1640
rect 415 1360 425 1630
rect 445 1360 455 1630
rect 415 1350 455 1360
rect 515 1630 555 1640
rect 515 1360 525 1630
rect 545 1360 555 1630
rect 515 1350 555 1360
rect 615 1630 655 1640
rect 615 1360 625 1630
rect 645 1360 655 1630
rect 615 1350 655 1360
rect 715 1630 755 1640
rect 715 1360 725 1630
rect 745 1360 755 1630
rect 715 1350 755 1360
rect 815 1630 855 1640
rect 815 1360 825 1630
rect 845 1360 855 1630
rect 815 1350 855 1360
rect 915 1630 955 1640
rect 915 1360 925 1630
rect 945 1360 955 1630
rect 915 1350 955 1360
rect 1015 1630 1055 1640
rect 1015 1360 1025 1630
rect 1045 1360 1055 1630
rect 1015 1350 1055 1360
rect 1115 1630 1155 1640
rect 1115 1360 1125 1630
rect 1145 1360 1155 1630
rect 1115 1350 1155 1360
rect 225 1135 245 1350
rect 425 1135 445 1350
rect 625 1135 645 1350
rect 825 1135 845 1350
rect 1025 1135 1045 1350
rect 115 1125 155 1135
rect 115 855 125 1125
rect 145 855 155 1125
rect 115 845 155 855
rect 215 1125 255 1135
rect 215 855 225 1125
rect 245 855 255 1125
rect 215 845 255 855
rect 315 1125 355 1135
rect 315 855 325 1125
rect 345 855 355 1125
rect 315 845 355 855
rect 415 1125 455 1135
rect 415 855 425 1125
rect 445 855 455 1125
rect 415 845 455 855
rect 515 1125 555 1135
rect 515 855 525 1125
rect 545 855 555 1125
rect 515 845 555 855
rect 615 1125 655 1135
rect 615 855 625 1125
rect 645 855 655 1125
rect 615 845 655 855
rect 715 1125 755 1135
rect 715 855 725 1125
rect 745 855 755 1125
rect 715 845 755 855
rect 815 1125 855 1135
rect 815 855 825 1125
rect 845 855 855 1125
rect 815 845 855 855
rect 915 1125 955 1135
rect 915 855 925 1125
rect 945 855 955 1125
rect 915 845 955 855
rect 1015 1125 1055 1135
rect 1015 855 1025 1125
rect 1045 855 1055 1125
rect 1015 845 1055 855
rect 1115 1125 1155 1135
rect 1115 855 1125 1125
rect 1145 855 1155 1125
rect 1115 845 1155 855
rect 165 815 205 825
rect 165 795 175 815
rect 195 795 205 815
rect 165 785 205 795
rect 5 740 45 750
rect 5 720 15 740
rect 35 720 45 740
rect 225 730 245 845
rect 425 730 445 845
rect 5 710 45 720
rect 65 710 245 730
rect 345 710 445 730
rect 65 690 85 710
rect 345 690 365 710
rect 625 690 645 845
rect 825 730 845 845
rect 1025 730 1045 845
rect 1065 815 1105 825
rect 1065 795 1075 815
rect 1095 795 1105 815
rect 1065 785 1105 795
rect 1225 740 1265 750
rect 825 710 925 730
rect 1025 710 1205 730
rect 1225 720 1235 740
rect 1255 720 1265 740
rect 1225 710 1265 720
rect 905 690 925 710
rect 1185 690 1205 710
rect -45 680 -5 690
rect -45 410 -35 680
rect -15 410 -5 680
rect -45 400 -5 410
rect 55 680 95 690
rect 55 410 65 680
rect 85 410 95 680
rect 55 400 95 410
rect 155 680 195 690
rect 155 410 165 680
rect 185 410 195 680
rect 155 400 195 410
rect 235 680 275 690
rect 235 410 245 680
rect 265 410 275 680
rect 235 400 275 410
rect 335 680 375 690
rect 335 410 345 680
rect 365 410 375 680
rect 335 400 375 410
rect 435 680 475 690
rect 435 410 445 680
rect 465 410 475 680
rect 435 400 475 410
rect 515 680 555 690
rect 515 410 525 680
rect 545 410 555 680
rect 515 400 555 410
rect 615 680 655 690
rect 615 410 625 680
rect 645 410 655 680
rect 615 400 655 410
rect 715 680 755 690
rect 715 410 725 680
rect 745 410 755 680
rect 715 400 755 410
rect 795 680 835 690
rect 795 410 805 680
rect 825 410 835 680
rect 795 400 835 410
rect 895 680 935 690
rect 895 410 905 680
rect 925 410 935 680
rect 895 400 935 410
rect 995 680 1035 690
rect 995 410 1005 680
rect 1025 410 1035 680
rect 995 400 1035 410
rect 1075 680 1115 690
rect 1075 410 1085 680
rect 1105 410 1115 680
rect 1075 400 1115 410
rect 1175 680 1215 690
rect 1175 410 1185 680
rect 1205 410 1215 680
rect 1175 400 1215 410
rect 1275 680 1315 690
rect 1275 410 1285 680
rect 1305 410 1315 680
rect 1275 400 1315 410
rect 175 335 195 400
rect 245 375 265 400
rect 455 375 475 400
rect 245 355 475 375
rect 245 335 265 355
rect 455 335 475 355
rect 535 375 555 400
rect 725 375 745 400
rect 535 355 745 375
rect 535 335 555 355
rect 725 335 745 355
rect 805 375 825 400
rect 1005 375 1025 400
rect 805 355 1025 375
rect 805 335 825 355
rect 1005 335 1025 355
rect 1075 335 1095 400
rect -45 325 -5 335
rect -45 55 -35 325
rect -15 55 -5 325
rect -45 45 -5 55
rect 55 325 95 335
rect 55 55 65 325
rect 85 55 95 325
rect 55 45 95 55
rect 155 325 195 335
rect 155 55 165 325
rect 185 55 195 325
rect 155 45 195 55
rect 235 325 275 335
rect 235 55 245 325
rect 265 55 275 325
rect 235 45 275 55
rect 335 325 375 335
rect 335 55 345 325
rect 365 55 375 325
rect 335 45 375 55
rect 435 325 475 335
rect 435 55 445 325
rect 465 55 475 325
rect 435 45 475 55
rect 515 325 555 335
rect 515 55 525 325
rect 545 55 555 325
rect 515 45 555 55
rect 615 325 655 335
rect 615 55 625 325
rect 645 55 655 325
rect 615 45 655 55
rect 715 325 755 335
rect 715 55 725 325
rect 745 55 755 325
rect 715 45 755 55
rect 795 325 835 335
rect 795 55 805 325
rect 825 55 835 325
rect 795 45 835 55
rect 895 325 935 335
rect 895 55 905 325
rect 925 55 935 325
rect 895 45 935 55
rect 995 325 1035 335
rect 995 55 1005 325
rect 1025 55 1035 325
rect 995 45 1035 55
rect 1075 325 1115 335
rect 1075 55 1085 325
rect 1105 55 1115 325
rect 1075 45 1115 55
rect 1175 325 1215 335
rect 1175 55 1185 325
rect 1205 55 1215 325
rect 1175 45 1215 55
rect 1275 325 1315 335
rect 1275 55 1285 325
rect 1305 55 1315 325
rect 1275 45 1315 55
rect 5 15 45 25
rect 5 -5 15 15
rect 35 -5 45 15
rect 105 15 145 25
rect 105 5 115 15
rect 5 -15 45 -5
rect 65 -5 115 5
rect 135 -5 145 15
rect 65 -15 145 -5
rect 1225 15 1265 25
rect 1225 -5 1235 15
rect 1255 -5 1265 15
rect 1225 -15 1265 -5
rect 65 -35 85 -15
rect 25 -55 85 -35
rect 115 -80 155 -70
rect 115 -350 125 -80
rect 145 -350 155 -80
rect 115 -360 155 -350
rect 215 -80 255 -70
rect 215 -350 225 -80
rect 245 -350 255 -80
rect 215 -360 255 -350
rect 315 -80 355 -70
rect 315 -350 325 -80
rect 345 -350 355 -80
rect 315 -360 355 -350
rect 415 -80 455 -70
rect 415 -350 425 -80
rect 445 -350 455 -80
rect 415 -360 455 -350
rect 515 -80 555 -70
rect 515 -350 525 -80
rect 545 -350 555 -80
rect 515 -360 555 -350
rect 615 -80 655 -70
rect 615 -350 625 -80
rect 645 -350 655 -80
rect 615 -360 655 -350
rect 715 -80 755 -70
rect 715 -350 725 -80
rect 745 -350 755 -80
rect 715 -360 755 -350
rect 815 -80 855 -70
rect 815 -350 825 -80
rect 845 -350 855 -80
rect 815 -360 855 -350
rect 915 -80 955 -70
rect 915 -350 925 -80
rect 945 -350 955 -80
rect 915 -360 955 -350
rect 1015 -80 1055 -70
rect 1015 -350 1025 -80
rect 1045 -350 1055 -80
rect 1015 -360 1055 -350
rect 1115 -80 1155 -70
rect 1115 -350 1125 -80
rect 1145 -350 1155 -80
rect 1115 -360 1155 -350
rect 165 -390 205 -380
rect 165 -410 175 -390
rect 195 -410 205 -390
rect 165 -420 205 -410
rect 1065 -390 1105 -380
rect 1065 -410 1075 -390
rect 1095 -410 1105 -390
rect 1065 -420 1105 -410
<< viali >>
rect 125 1795 145 2065
rect 325 1795 345 2065
rect 525 1795 545 2065
rect 725 1795 745 2065
rect 925 1795 945 2065
rect 1125 1795 1145 2065
rect 125 1360 145 1630
rect 225 1360 245 1380
rect 425 1390 445 1410
rect 625 1360 645 1380
rect 825 1390 845 1410
rect 1025 1360 1045 1380
rect 1125 1360 1145 1630
rect 125 855 145 1125
rect 325 855 345 1125
rect 525 855 545 1125
rect 725 855 745 1125
rect 925 855 945 1125
rect 1125 855 1145 1125
rect 65 305 85 325
rect 165 245 185 265
rect 345 275 365 295
rect 445 190 465 210
rect 525 220 545 240
rect 625 305 645 325
rect 725 220 745 240
rect 805 190 825 210
rect 905 275 925 295
rect 1085 245 1105 265
rect 1185 305 1205 325
rect 125 -350 145 -80
rect 325 -350 345 -80
rect 525 -350 545 -80
rect 725 -350 745 -80
rect 925 -350 945 -80
rect 1125 -350 1145 -80
<< metal1 >>
rect 415 1410 855 1420
rect 415 1390 425 1410
rect 445 1405 825 1410
rect 445 1390 455 1405
rect 815 1390 825 1405
rect 845 1390 855 1410
rect 215 1380 255 1390
rect 415 1380 455 1390
rect 615 1380 655 1390
rect 815 1380 855 1390
rect 1015 1380 1055 1390
rect 215 1360 225 1380
rect 245 1365 255 1380
rect 615 1365 625 1380
rect 245 1360 625 1365
rect 645 1365 655 1380
rect 1015 1365 1025 1380
rect 645 1360 1025 1365
rect 1045 1360 1055 1380
rect 215 1350 1055 1360
rect 55 325 1215 335
rect 55 305 65 325
rect 85 320 625 325
rect 85 305 95 320
rect 615 305 625 320
rect 645 320 1185 325
rect 645 305 655 320
rect 1175 305 1185 320
rect 1205 305 1215 325
rect 55 295 95 305
rect 335 295 375 305
rect 615 295 655 305
rect 895 295 935 305
rect 1175 295 1215 305
rect 335 275 345 295
rect 365 280 375 295
rect 895 280 905 295
rect 365 275 905 280
rect 925 275 935 295
rect 155 265 195 275
rect 335 265 935 275
rect 1075 265 1115 275
rect 155 245 165 265
rect 185 250 195 265
rect 1075 250 1085 265
rect 185 245 1085 250
rect 1105 245 1115 265
rect 155 240 1115 245
rect 155 235 525 240
rect 515 220 525 235
rect 545 235 725 240
rect 545 220 555 235
rect 435 210 475 220
rect 515 210 555 220
rect 715 220 725 235
rect 745 235 1115 240
rect 745 220 755 235
rect 715 210 755 220
rect 795 210 835 220
rect 435 190 445 210
rect 465 195 475 210
rect 795 195 805 210
rect 465 190 805 195
rect 825 190 835 210
rect 435 180 835 190
<< end >>
