* SPICE3 file created from shiftregister_inverter.ext - technology: sky130A

.subckt shiftregister_inverter VP
X0 a_n160_730# a_n420_730# a_n290_730# VSUBS sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X1 a_n160_730# a_n420_730# a_n290_1070# VP sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=0.5 ps=2.5 w=2 l=0.15
X2 a_n290_730# A a_n420_730# VSUBS sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.15
X3 a_n290_1070# A a_n420_1070# VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=1 ps=5 w=2 l=0.15
.ends
