magic
tech sky130A
timestamp 1697145733
<< error_p >>
rect -325 1552 -65 1555
rect -325 1288 -322 1552
rect -68 1288 -65 1552
rect -325 1285 -65 1288
rect 1815 1552 2075 1555
rect 1815 1288 1818 1552
rect 2072 1288 2075 1552
rect 1815 1285 2075 1288
rect -125 1102 -105 1105
rect -125 838 -122 1102
rect -108 838 -105 1102
rect -125 835 -105 838
rect 75 1102 95 1105
rect 75 838 78 1102
rect 92 838 95 1102
rect 75 835 95 838
rect 255 1102 275 1105
rect 255 838 258 1102
rect 272 838 275 1102
rect 255 835 275 838
rect 305 1102 325 1105
rect 305 838 308 1102
rect 322 838 325 1102
rect 305 835 325 838
rect 865 1102 885 1105
rect 865 838 868 1102
rect 882 838 885 1102
rect 865 835 885 838
rect 1245 1102 1265 1105
rect 1245 838 1248 1102
rect 1262 838 1265 1102
rect 1245 835 1265 838
rect 1425 1102 1445 1105
rect 1425 838 1428 1102
rect 1442 838 1445 1102
rect 1425 835 1445 838
rect 1475 1102 1495 1105
rect 1475 838 1478 1102
rect 1492 838 1495 1102
rect 1475 835 1495 838
rect -125 712 -105 715
rect -125 448 -122 712
rect -108 448 -105 712
rect -125 445 -105 448
rect 75 712 95 715
rect 75 448 78 712
rect 92 448 95 712
rect 75 445 95 448
rect 255 712 275 715
rect 255 448 258 712
rect 272 448 275 712
rect 255 445 275 448
rect 305 712 325 715
rect 305 448 308 712
rect 322 448 325 712
rect 305 445 325 448
rect 865 712 885 715
rect 865 448 868 712
rect 882 448 885 712
rect 865 445 885 448
rect 1245 712 1265 715
rect 1245 448 1248 712
rect 1262 448 1265 712
rect 1245 445 1265 448
rect 1425 712 1445 715
rect 1425 448 1428 712
rect 1442 448 1445 712
rect 1425 445 1445 448
rect 1475 712 1495 715
rect 1475 448 1478 712
rect 1492 448 1495 712
rect 1475 445 1495 448
rect -325 262 -65 265
rect -325 -2 -322 262
rect -68 -2 -65 262
rect -325 -5 -65 -2
rect 1815 262 2075 265
rect 1815 -2 1818 262
rect 2072 -2 2075 262
rect 1815 -5 2075 -2
<< nwell >>
rect -360 800 2110 1590
<< nmos >>
rect -290 430 -240 730
rect -190 430 -140 730
rect -90 430 -40 730
rect 10 430 60 730
rect 110 430 160 730
rect 340 430 390 730
rect 520 430 570 730
rect 620 430 670 730
rect 800 430 850 730
rect 900 430 950 730
rect 1080 430 1130 730
rect 1180 430 1230 730
rect 1360 430 1410 730
rect 1590 430 1640 730
rect 1690 430 1740 730
rect 1790 430 1840 730
rect 1890 430 1940 730
rect 1990 430 2040 730
rect 0 -20 50 280
rect 100 -20 150 280
rect 200 -20 250 280
rect 300 -20 350 280
rect 400 -20 450 280
rect 500 -20 550 280
rect 600 -20 650 280
rect 700 -20 750 280
rect 800 -20 850 280
rect 900 -20 950 280
rect 1000 -20 1050 280
rect 1100 -20 1150 280
rect 1200 -20 1250 280
rect 1300 -20 1350 280
rect 1400 -20 1450 280
rect 1500 -20 1550 280
rect 1600 -20 1650 280
rect 1700 -20 1750 280
<< pmos >>
rect 0 1270 50 1570
rect 100 1270 150 1570
rect 200 1270 250 1570
rect 300 1270 350 1570
rect 400 1270 450 1570
rect 500 1270 550 1570
rect 600 1270 650 1570
rect 700 1270 750 1570
rect 800 1270 850 1570
rect 900 1270 950 1570
rect 1000 1270 1050 1570
rect 1100 1270 1150 1570
rect 1200 1270 1250 1570
rect 1300 1270 1350 1570
rect 1400 1270 1450 1570
rect 1500 1270 1550 1570
rect 1600 1270 1650 1570
rect 1700 1270 1750 1570
rect -290 820 -240 1120
rect -190 820 -140 1120
rect -90 820 -40 1120
rect 10 820 60 1120
rect 110 820 160 1120
rect 340 820 390 1120
rect 520 820 570 1120
rect 620 820 670 1120
rect 800 820 850 1120
rect 900 820 950 1120
rect 1080 820 1130 1120
rect 1180 820 1230 1120
rect 1360 820 1410 1120
rect 1590 820 1640 1120
rect 1690 820 1740 1120
rect 1790 820 1840 1120
rect 1890 820 1940 1120
rect 1990 820 2040 1120
<< ndiff >>
rect -340 715 -290 730
rect -340 445 -325 715
rect -305 445 -290 715
rect -340 430 -290 445
rect -240 715 -190 730
rect -240 445 -225 715
rect -205 445 -190 715
rect -240 430 -190 445
rect -140 715 -90 730
rect -140 445 -125 715
rect -105 445 -90 715
rect -140 430 -90 445
rect -40 715 10 730
rect -40 445 -25 715
rect -5 445 10 715
rect -40 430 10 445
rect 60 715 110 730
rect 60 445 75 715
rect 95 445 110 715
rect 60 430 110 445
rect 160 715 210 730
rect 160 445 175 715
rect 195 445 210 715
rect 160 430 210 445
rect 290 715 340 730
rect 290 445 305 715
rect 325 445 340 715
rect 290 430 340 445
rect 390 715 440 730
rect 390 445 405 715
rect 425 445 440 715
rect 390 430 440 445
rect 470 715 520 730
rect 470 445 485 715
rect 505 445 520 715
rect 470 430 520 445
rect 570 715 620 730
rect 570 445 585 715
rect 605 445 620 715
rect 570 430 620 445
rect 670 715 720 730
rect 670 445 685 715
rect 705 445 720 715
rect 670 430 720 445
rect 750 715 800 730
rect 750 445 765 715
rect 785 445 800 715
rect 750 430 800 445
rect 850 715 900 730
rect 850 445 865 715
rect 885 445 900 715
rect 850 430 900 445
rect 950 715 1000 730
rect 950 445 965 715
rect 985 445 1000 715
rect 950 430 1000 445
rect 1030 715 1080 730
rect 1030 445 1045 715
rect 1065 445 1080 715
rect 1030 430 1080 445
rect 1130 715 1180 730
rect 1130 445 1145 715
rect 1165 445 1180 715
rect 1130 430 1180 445
rect 1230 715 1280 730
rect 1230 445 1245 715
rect 1265 445 1280 715
rect 1230 430 1280 445
rect 1310 715 1360 730
rect 1310 445 1325 715
rect 1345 445 1360 715
rect 1310 430 1360 445
rect 1410 715 1460 730
rect 1410 445 1425 715
rect 1445 445 1460 715
rect 1410 430 1460 445
rect 1540 715 1590 730
rect 1540 445 1555 715
rect 1575 445 1590 715
rect 1540 430 1590 445
rect 1640 715 1690 730
rect 1640 445 1655 715
rect 1675 445 1690 715
rect 1640 430 1690 445
rect 1740 715 1790 730
rect 1740 445 1755 715
rect 1775 445 1790 715
rect 1740 430 1790 445
rect 1840 715 1890 730
rect 1840 445 1855 715
rect 1875 445 1890 715
rect 1840 430 1890 445
rect 1940 715 1990 730
rect 1940 445 1955 715
rect 1975 445 1990 715
rect 1940 430 1990 445
rect 2040 715 2090 730
rect 2040 445 2055 715
rect 2075 445 2090 715
rect 2040 430 2090 445
rect -50 265 0 280
rect -50 -5 -35 265
rect -15 -5 0 265
rect -50 -20 0 -5
rect 50 265 100 280
rect 50 -5 65 265
rect 85 -5 100 265
rect 50 -20 100 -5
rect 150 265 200 280
rect 150 -5 165 265
rect 185 -5 200 265
rect 150 -20 200 -5
rect 250 265 300 280
rect 250 -5 265 265
rect 285 -5 300 265
rect 250 -20 300 -5
rect 350 265 400 280
rect 350 -5 365 265
rect 385 -5 400 265
rect 350 -20 400 -5
rect 450 265 500 280
rect 450 -5 465 265
rect 485 -5 500 265
rect 450 -20 500 -5
rect 550 265 600 280
rect 550 -5 565 265
rect 585 -5 600 265
rect 550 -20 600 -5
rect 650 265 700 280
rect 650 -5 665 265
rect 685 -5 700 265
rect 650 -20 700 -5
rect 750 265 800 280
rect 750 -5 765 265
rect 785 -5 800 265
rect 750 -20 800 -5
rect 850 265 900 280
rect 850 -5 865 265
rect 885 -5 900 265
rect 850 -20 900 -5
rect 950 265 1000 280
rect 950 -5 965 265
rect 985 -5 1000 265
rect 950 -20 1000 -5
rect 1050 265 1100 280
rect 1050 -5 1065 265
rect 1085 -5 1100 265
rect 1050 -20 1100 -5
rect 1150 265 1200 280
rect 1150 -5 1165 265
rect 1185 -5 1200 265
rect 1150 -20 1200 -5
rect 1250 265 1300 280
rect 1250 -5 1265 265
rect 1285 -5 1300 265
rect 1250 -20 1300 -5
rect 1350 265 1400 280
rect 1350 -5 1365 265
rect 1385 -5 1400 265
rect 1350 -20 1400 -5
rect 1450 265 1500 280
rect 1450 -5 1465 265
rect 1485 -5 1500 265
rect 1450 -20 1500 -5
rect 1550 265 1600 280
rect 1550 -5 1565 265
rect 1585 -5 1600 265
rect 1550 -20 1600 -5
rect 1650 265 1700 280
rect 1650 -5 1665 265
rect 1685 -5 1700 265
rect 1650 -20 1700 -5
rect 1750 265 1800 280
rect 1750 -5 1765 265
rect 1785 -5 1800 265
rect 1750 -20 1800 -5
<< pdiff >>
rect -50 1555 0 1570
rect -50 1285 -35 1555
rect -15 1285 0 1555
rect -50 1270 0 1285
rect 50 1555 100 1570
rect 50 1285 65 1555
rect 85 1285 100 1555
rect 50 1270 100 1285
rect 150 1555 200 1570
rect 150 1285 165 1555
rect 185 1285 200 1555
rect 150 1270 200 1285
rect 250 1555 300 1570
rect 250 1285 265 1555
rect 285 1285 300 1555
rect 250 1270 300 1285
rect 350 1555 400 1570
rect 350 1285 365 1555
rect 385 1285 400 1555
rect 350 1270 400 1285
rect 450 1555 500 1570
rect 450 1285 465 1555
rect 485 1285 500 1555
rect 450 1270 500 1285
rect 550 1555 600 1570
rect 550 1285 565 1555
rect 585 1285 600 1555
rect 550 1270 600 1285
rect 650 1555 700 1570
rect 650 1285 665 1555
rect 685 1285 700 1555
rect 650 1270 700 1285
rect 750 1555 800 1570
rect 750 1285 765 1555
rect 785 1285 800 1555
rect 750 1270 800 1285
rect 850 1555 900 1570
rect 850 1285 865 1555
rect 885 1285 900 1555
rect 850 1270 900 1285
rect 950 1555 1000 1570
rect 950 1285 965 1555
rect 985 1285 1000 1555
rect 950 1270 1000 1285
rect 1050 1555 1100 1570
rect 1050 1285 1065 1555
rect 1085 1285 1100 1555
rect 1050 1270 1100 1285
rect 1150 1555 1200 1570
rect 1150 1285 1165 1555
rect 1185 1285 1200 1555
rect 1150 1270 1200 1285
rect 1250 1555 1300 1570
rect 1250 1285 1265 1555
rect 1285 1285 1300 1555
rect 1250 1270 1300 1285
rect 1350 1555 1400 1570
rect 1350 1285 1365 1555
rect 1385 1285 1400 1555
rect 1350 1270 1400 1285
rect 1450 1555 1500 1570
rect 1450 1285 1465 1555
rect 1485 1285 1500 1555
rect 1450 1270 1500 1285
rect 1550 1555 1600 1570
rect 1550 1285 1565 1555
rect 1585 1285 1600 1555
rect 1550 1270 1600 1285
rect 1650 1555 1700 1570
rect 1650 1285 1665 1555
rect 1685 1285 1700 1555
rect 1650 1270 1700 1285
rect 1750 1555 1800 1570
rect 1750 1285 1765 1555
rect 1785 1285 1800 1555
rect 1750 1270 1800 1285
rect -340 1105 -290 1120
rect -340 835 -325 1105
rect -305 835 -290 1105
rect -340 820 -290 835
rect -240 1105 -190 1120
rect -240 835 -225 1105
rect -205 835 -190 1105
rect -240 820 -190 835
rect -140 1105 -90 1120
rect -140 835 -125 1105
rect -105 835 -90 1105
rect -140 820 -90 835
rect -40 1105 10 1120
rect -40 835 -25 1105
rect -5 835 10 1105
rect -40 820 10 835
rect 60 1105 110 1120
rect 60 835 75 1105
rect 95 835 110 1105
rect 60 820 110 835
rect 160 1105 210 1120
rect 160 835 175 1105
rect 195 835 210 1105
rect 160 820 210 835
rect 290 1105 340 1120
rect 290 835 305 1105
rect 325 835 340 1105
rect 290 820 340 835
rect 390 1105 440 1120
rect 390 835 405 1105
rect 425 835 440 1105
rect 390 820 440 835
rect 470 1105 520 1120
rect 470 835 485 1105
rect 505 835 520 1105
rect 470 820 520 835
rect 570 1105 620 1120
rect 570 835 585 1105
rect 605 835 620 1105
rect 570 820 620 835
rect 670 1105 720 1120
rect 670 835 685 1105
rect 705 835 720 1105
rect 670 820 720 835
rect 750 1105 800 1120
rect 750 835 765 1105
rect 785 835 800 1105
rect 750 820 800 835
rect 850 1105 900 1120
rect 850 835 865 1105
rect 885 835 900 1105
rect 850 820 900 835
rect 950 1105 1000 1120
rect 950 835 965 1105
rect 985 835 1000 1105
rect 950 820 1000 835
rect 1030 1105 1080 1120
rect 1030 835 1045 1105
rect 1065 835 1080 1105
rect 1030 820 1080 835
rect 1130 1105 1180 1120
rect 1130 835 1145 1105
rect 1165 835 1180 1105
rect 1130 820 1180 835
rect 1230 1105 1280 1120
rect 1230 835 1245 1105
rect 1265 835 1280 1105
rect 1230 820 1280 835
rect 1310 1105 1360 1120
rect 1310 835 1325 1105
rect 1345 835 1360 1105
rect 1310 820 1360 835
rect 1410 1105 1460 1120
rect 1410 835 1425 1105
rect 1445 835 1460 1105
rect 1410 820 1460 835
rect 1540 1105 1590 1120
rect 1540 835 1555 1105
rect 1575 835 1590 1105
rect 1540 820 1590 835
rect 1640 1105 1690 1120
rect 1640 835 1655 1105
rect 1675 835 1690 1105
rect 1640 820 1690 835
rect 1740 1105 1790 1120
rect 1740 835 1755 1105
rect 1775 835 1790 1105
rect 1740 820 1790 835
rect 1840 1105 1890 1120
rect 1840 835 1855 1105
rect 1875 835 1890 1105
rect 1840 820 1890 835
rect 1940 1105 1990 1120
rect 1940 835 1955 1105
rect 1975 835 1990 1105
rect 1940 820 1990 835
rect 2040 1105 2090 1120
rect 2040 835 2055 1105
rect 2075 835 2090 1105
rect 2040 820 2090 835
<< ndiffc >>
rect -325 445 -305 715
rect -225 445 -205 715
rect -125 445 -105 715
rect -25 445 -5 715
rect 75 445 95 715
rect 175 445 195 715
rect 305 445 325 715
rect 405 445 425 715
rect 485 445 505 715
rect 585 445 605 715
rect 685 445 705 715
rect 765 445 785 715
rect 865 445 885 715
rect 965 445 985 715
rect 1045 445 1065 715
rect 1145 445 1165 715
rect 1245 445 1265 715
rect 1325 445 1345 715
rect 1425 445 1445 715
rect 1555 445 1575 715
rect 1655 445 1675 715
rect 1755 445 1775 715
rect 1855 445 1875 715
rect 1955 445 1975 715
rect 2055 445 2075 715
rect -35 -5 -15 265
rect 65 -5 85 265
rect 165 -5 185 265
rect 265 -5 285 265
rect 365 -5 385 265
rect 465 -5 485 265
rect 565 -5 585 265
rect 665 -5 685 265
rect 765 -5 785 265
rect 865 -5 885 265
rect 965 -5 985 265
rect 1065 -5 1085 265
rect 1165 -5 1185 265
rect 1265 -5 1285 265
rect 1365 -5 1385 265
rect 1465 -5 1485 265
rect 1565 -5 1585 265
rect 1665 -5 1685 265
rect 1765 -5 1785 265
<< pdiffc >>
rect -35 1285 -15 1555
rect 65 1285 85 1555
rect 165 1285 185 1555
rect 265 1285 285 1555
rect 365 1285 385 1555
rect 465 1285 485 1555
rect 565 1285 585 1555
rect 665 1285 685 1555
rect 765 1285 785 1555
rect 865 1285 885 1555
rect 965 1285 985 1555
rect 1065 1285 1085 1555
rect 1165 1285 1185 1555
rect 1265 1285 1285 1555
rect 1365 1285 1385 1555
rect 1465 1285 1485 1555
rect 1565 1285 1585 1555
rect 1665 1285 1685 1555
rect 1765 1285 1785 1555
rect -325 835 -305 1105
rect -225 835 -205 1105
rect -125 835 -105 1105
rect -25 835 -5 1105
rect 75 835 95 1105
rect 175 835 195 1105
rect 305 835 325 1105
rect 405 835 425 1105
rect 485 835 505 1105
rect 585 835 605 1105
rect 685 835 705 1105
rect 765 835 785 1105
rect 865 835 885 1105
rect 965 835 985 1105
rect 1045 835 1065 1105
rect 1145 835 1165 1105
rect 1245 835 1265 1105
rect 1325 835 1345 1105
rect 1425 835 1445 1105
rect 1555 835 1575 1105
rect 1655 835 1675 1105
rect 1755 835 1775 1105
rect 1855 835 1875 1105
rect 1955 835 1975 1105
rect 2055 835 2075 1105
<< psubdiff >>
rect 240 715 290 730
rect 240 445 255 715
rect 275 445 290 715
rect 240 430 290 445
rect 1460 715 1510 730
rect 1460 445 1475 715
rect 1495 445 1510 715
rect 1460 430 1510 445
rect -340 265 -50 280
rect -340 -5 -325 265
rect -65 -5 -50 265
rect -340 -20 -50 -5
rect 1800 265 2090 280
rect 1800 -5 1815 265
rect 2075 -5 2090 265
rect 1800 -20 2090 -5
<< nsubdiff >>
rect -340 1555 -50 1570
rect -340 1285 -325 1555
rect -65 1285 -50 1555
rect -340 1270 -50 1285
rect 1800 1555 2090 1570
rect 1800 1285 1815 1555
rect 2075 1285 2090 1555
rect 1800 1270 2090 1285
rect 240 1105 290 1120
rect 240 835 255 1105
rect 275 835 290 1105
rect 240 820 290 835
rect 1460 1105 1510 1120
rect 1460 835 1475 1105
rect 1495 835 1510 1105
rect 1460 820 1510 835
<< psubdiffcont >>
rect 255 445 275 715
rect 1475 445 1495 715
rect -325 -5 -65 265
rect 1815 -5 2075 265
<< nsubdiffcont >>
rect -325 1285 -65 1555
rect 1815 1285 2075 1555
rect 255 835 275 1105
rect 1475 835 1495 1105
<< poly >>
rect 0 1570 50 1585
rect 100 1570 150 1585
rect 200 1570 250 1585
rect 300 1570 350 1585
rect 400 1570 450 1585
rect 500 1570 550 1585
rect 600 1570 650 1585
rect 700 1570 750 1585
rect 800 1570 850 1585
rect 900 1570 950 1585
rect 1000 1570 1050 1585
rect 1100 1570 1150 1585
rect 1200 1570 1250 1585
rect 1300 1570 1350 1585
rect 1400 1570 1450 1585
rect 1500 1570 1550 1585
rect 1600 1570 1650 1585
rect 1700 1570 1750 1585
rect 0 1245 50 1270
rect 0 1225 15 1245
rect 35 1225 50 1245
rect 0 1215 50 1225
rect 100 1245 150 1270
rect 100 1225 115 1245
rect 135 1225 150 1245
rect 100 1215 150 1225
rect 200 1245 250 1270
rect 200 1225 215 1245
rect 235 1225 250 1245
rect 200 1215 250 1225
rect 300 1245 350 1270
rect 300 1225 315 1245
rect 335 1225 350 1245
rect 300 1215 350 1225
rect 400 1245 450 1270
rect 400 1225 415 1245
rect 435 1225 450 1245
rect 400 1215 450 1225
rect 500 1245 550 1270
rect 500 1225 515 1245
rect 535 1225 550 1245
rect 500 1215 550 1225
rect 600 1245 650 1270
rect 600 1225 615 1245
rect 635 1225 650 1245
rect 600 1215 650 1225
rect 700 1245 750 1270
rect 700 1225 715 1245
rect 735 1225 750 1245
rect 700 1215 750 1225
rect 800 1245 850 1270
rect 800 1225 815 1245
rect 835 1225 850 1245
rect 800 1215 850 1225
rect 900 1245 950 1270
rect 900 1225 915 1245
rect 935 1225 950 1245
rect 900 1215 950 1225
rect 1000 1245 1050 1270
rect 1000 1225 1015 1245
rect 1035 1225 1050 1245
rect 1000 1215 1050 1225
rect 1100 1245 1150 1270
rect 1100 1225 1115 1245
rect 1135 1225 1150 1245
rect 1100 1215 1150 1225
rect 1200 1245 1250 1270
rect 1200 1225 1215 1245
rect 1235 1225 1250 1245
rect 1200 1215 1250 1225
rect 1300 1245 1350 1270
rect 1300 1225 1315 1245
rect 1335 1225 1350 1245
rect 1300 1215 1350 1225
rect 1400 1245 1450 1270
rect 1400 1225 1415 1245
rect 1435 1225 1450 1245
rect 1400 1215 1450 1225
rect 1500 1245 1550 1270
rect 1500 1225 1515 1245
rect 1535 1225 1550 1245
rect 1500 1215 1550 1225
rect 1600 1245 1650 1270
rect 1600 1225 1615 1245
rect 1635 1225 1650 1245
rect 1600 1215 1650 1225
rect 1700 1245 1750 1270
rect 1700 1225 1715 1245
rect 1735 1225 1750 1245
rect 1700 1215 1750 1225
rect -290 1165 -240 1175
rect -290 1145 -275 1165
rect -255 1145 -240 1165
rect -290 1120 -240 1145
rect -190 1165 -140 1175
rect -190 1145 -175 1165
rect -155 1145 -140 1165
rect -190 1120 -140 1145
rect -90 1165 -40 1175
rect -90 1145 -75 1165
rect -55 1145 -40 1165
rect -90 1120 -40 1145
rect 10 1165 60 1175
rect 10 1145 25 1165
rect 45 1145 60 1165
rect 10 1120 60 1145
rect 110 1165 160 1175
rect 110 1145 125 1165
rect 145 1145 160 1165
rect 110 1120 160 1145
rect 340 1165 1410 1175
rect 340 1145 355 1165
rect 375 1145 1410 1165
rect 340 1135 1410 1145
rect 340 1120 390 1135
rect 520 1120 570 1135
rect 620 1120 670 1135
rect 800 1120 850 1135
rect 900 1120 950 1135
rect 1080 1120 1130 1135
rect 1180 1120 1230 1135
rect 1360 1120 1410 1135
rect 1590 1165 1640 1175
rect 1590 1145 1605 1165
rect 1625 1145 1640 1165
rect 1590 1120 1640 1145
rect 1690 1165 1740 1175
rect 1690 1145 1705 1165
rect 1725 1145 1740 1165
rect 1690 1120 1740 1145
rect 1790 1165 1840 1175
rect 1790 1145 1805 1165
rect 1825 1145 1840 1165
rect 1790 1120 1840 1145
rect 1890 1165 1940 1175
rect 1890 1145 1905 1165
rect 1925 1145 1940 1165
rect 1890 1120 1940 1145
rect 1990 1165 2040 1175
rect 1990 1145 2005 1165
rect 2025 1145 2040 1165
rect 1990 1120 2040 1145
rect -290 805 -240 820
rect -190 805 -140 820
rect -90 805 -40 820
rect 10 805 60 820
rect 110 805 160 820
rect 340 805 390 820
rect 520 805 570 820
rect 620 805 670 820
rect 800 805 850 820
rect 900 805 950 820
rect 1080 805 1130 820
rect 1180 805 1230 820
rect 1360 805 1410 820
rect 1590 805 1640 820
rect 1690 805 1740 820
rect 1790 805 1840 820
rect 1890 805 1940 820
rect 1990 805 2040 820
rect -290 730 -240 745
rect -190 730 -140 745
rect -90 730 -40 745
rect 10 730 60 745
rect 110 730 160 745
rect 340 730 390 745
rect 520 730 570 745
rect 620 730 670 745
rect 800 730 850 745
rect 900 730 950 745
rect 1080 730 1130 745
rect 1180 730 1230 745
rect 1360 730 1410 745
rect 1590 730 1640 745
rect 1690 730 1740 745
rect 1790 730 1840 745
rect 1890 730 1940 745
rect 1990 730 2040 745
rect -290 405 -240 430
rect -290 385 -275 405
rect -255 385 -240 405
rect -290 375 -240 385
rect -190 405 -140 430
rect -190 385 -175 405
rect -155 385 -140 405
rect -190 375 -140 385
rect -90 405 -40 430
rect -90 385 -75 405
rect -55 385 -40 405
rect -90 375 -40 385
rect 10 405 60 430
rect 10 385 25 405
rect 45 385 60 405
rect 10 375 60 385
rect 110 405 160 430
rect 110 385 125 405
rect 145 385 160 405
rect 110 375 160 385
rect 340 415 390 430
rect 520 415 570 430
rect 620 415 670 430
rect 800 415 850 430
rect 900 415 950 430
rect 1080 415 1130 430
rect 1180 415 1230 430
rect 1360 415 1410 430
rect 340 405 1410 415
rect 340 385 355 405
rect 375 385 1410 405
rect 340 375 1410 385
rect 1590 405 1640 430
rect 1590 385 1605 405
rect 1625 385 1640 405
rect 1590 375 1640 385
rect 1690 405 1740 430
rect 1690 385 1705 405
rect 1725 385 1740 405
rect 1690 375 1740 385
rect 1790 405 1840 430
rect 1790 385 1805 405
rect 1825 385 1840 405
rect 1790 375 1840 385
rect 1890 405 1940 430
rect 1890 385 1905 405
rect 1925 385 1940 405
rect 1890 375 1940 385
rect 1990 405 2040 430
rect 1990 385 2005 405
rect 2025 385 2040 405
rect 1990 375 2040 385
rect 0 325 50 335
rect 0 305 15 325
rect 35 305 50 325
rect 0 280 50 305
rect 100 325 150 335
rect 100 305 115 325
rect 135 305 150 325
rect 100 280 150 305
rect 200 325 250 335
rect 200 305 215 325
rect 235 305 250 325
rect 200 280 250 305
rect 300 325 350 335
rect 300 305 315 325
rect 335 305 350 325
rect 300 280 350 305
rect 400 325 450 335
rect 400 305 415 325
rect 435 305 450 325
rect 400 280 450 305
rect 500 325 550 335
rect 500 305 515 325
rect 535 305 550 325
rect 500 280 550 305
rect 600 325 650 335
rect 600 305 615 325
rect 635 305 650 325
rect 600 280 650 305
rect 700 325 750 335
rect 700 305 715 325
rect 735 305 750 325
rect 700 280 750 305
rect 800 325 850 335
rect 800 305 815 325
rect 835 305 850 325
rect 800 280 850 305
rect 900 325 950 335
rect 900 305 915 325
rect 935 305 950 325
rect 900 280 950 305
rect 1000 325 1050 335
rect 1000 305 1015 325
rect 1035 305 1050 325
rect 1000 280 1050 305
rect 1100 325 1150 335
rect 1100 305 1115 325
rect 1135 305 1150 325
rect 1100 280 1150 305
rect 1200 325 1250 335
rect 1200 305 1215 325
rect 1235 305 1250 325
rect 1200 280 1250 305
rect 1300 325 1350 335
rect 1300 305 1315 325
rect 1335 305 1350 325
rect 1300 280 1350 305
rect 1400 325 1450 335
rect 1400 305 1415 325
rect 1435 305 1450 325
rect 1400 280 1450 305
rect 1500 325 1550 335
rect 1500 305 1515 325
rect 1535 305 1550 325
rect 1500 280 1550 305
rect 1600 325 1650 335
rect 1600 305 1615 325
rect 1635 305 1650 325
rect 1600 280 1650 305
rect 1700 325 1750 335
rect 1700 305 1715 325
rect 1735 305 1750 325
rect 1700 280 1750 305
rect 0 -35 50 -20
rect 100 -35 150 -20
rect 200 -35 250 -20
rect 300 -35 350 -20
rect 400 -35 450 -20
rect 500 -35 550 -20
rect 600 -35 650 -20
rect 700 -35 750 -20
rect 800 -35 850 -20
rect 900 -35 950 -20
rect 1000 -35 1050 -20
rect 1100 -35 1150 -20
rect 1200 -35 1250 -20
rect 1300 -35 1350 -20
rect 1400 -35 1450 -20
rect 1500 -35 1550 -20
rect 1600 -35 1650 -20
rect 1700 -35 1750 -20
<< polycont >>
rect 15 1225 35 1245
rect 115 1225 135 1245
rect 215 1225 235 1245
rect 315 1225 335 1245
rect 415 1225 435 1245
rect 515 1225 535 1245
rect 615 1225 635 1245
rect 715 1225 735 1245
rect 815 1225 835 1245
rect 915 1225 935 1245
rect 1015 1225 1035 1245
rect 1115 1225 1135 1245
rect 1215 1225 1235 1245
rect 1315 1225 1335 1245
rect 1415 1225 1435 1245
rect 1515 1225 1535 1245
rect 1615 1225 1635 1245
rect 1715 1225 1735 1245
rect -275 1145 -255 1165
rect -175 1145 -155 1165
rect -75 1145 -55 1165
rect 25 1145 45 1165
rect 125 1145 145 1165
rect 355 1145 375 1165
rect 1605 1145 1625 1165
rect 1705 1145 1725 1165
rect 1805 1145 1825 1165
rect 1905 1145 1925 1165
rect 2005 1145 2025 1165
rect -275 385 -255 405
rect -175 385 -155 405
rect -75 385 -55 405
rect 25 385 45 405
rect 125 385 145 405
rect 355 385 375 405
rect 1605 385 1625 405
rect 1705 385 1725 405
rect 1805 385 1825 405
rect 1905 385 1925 405
rect 2005 385 2025 405
rect 15 305 35 325
rect 115 305 135 325
rect 215 305 235 325
rect 315 305 335 325
rect 415 305 435 325
rect 515 305 535 325
rect 615 305 635 325
rect 715 305 735 325
rect 815 305 835 325
rect 915 305 935 325
rect 1015 305 1035 325
rect 1115 305 1135 325
rect 1215 305 1235 325
rect 1315 305 1335 325
rect 1415 305 1435 325
rect 1515 305 1535 325
rect 1615 305 1635 325
rect 1715 305 1735 325
<< locali >>
rect 65 1585 1685 1605
rect 65 1565 85 1585
rect 265 1565 285 1585
rect 465 1565 485 1585
rect 665 1565 685 1585
rect 865 1565 885 1585
rect 1065 1565 1085 1585
rect 1265 1565 1285 1585
rect 1465 1565 1485 1585
rect 1665 1565 1685 1585
rect -335 1555 -5 1565
rect -335 1285 -325 1555
rect -65 1285 -35 1555
rect -15 1285 -5 1555
rect -335 1275 -5 1285
rect 55 1555 95 1565
rect 55 1285 65 1555
rect 85 1285 95 1555
rect 55 1275 95 1285
rect 155 1555 195 1565
rect 155 1285 165 1555
rect 185 1285 195 1555
rect 155 1275 195 1285
rect 255 1555 295 1565
rect 255 1285 265 1555
rect 285 1285 295 1555
rect 255 1275 295 1285
rect 355 1555 395 1565
rect 355 1285 365 1555
rect 385 1285 395 1555
rect 355 1275 395 1285
rect 455 1555 495 1565
rect 455 1285 465 1555
rect 485 1285 495 1555
rect 455 1275 495 1285
rect 555 1555 595 1565
rect 555 1285 565 1555
rect 585 1285 595 1555
rect 555 1275 595 1285
rect 655 1555 695 1565
rect 655 1285 665 1555
rect 685 1285 695 1555
rect 655 1275 695 1285
rect 755 1555 795 1565
rect 755 1285 765 1555
rect 785 1285 795 1555
rect 755 1275 795 1285
rect 855 1555 895 1565
rect 855 1285 865 1555
rect 885 1285 895 1555
rect 855 1275 895 1285
rect 955 1555 995 1565
rect 955 1285 965 1555
rect 985 1285 995 1555
rect 955 1275 995 1285
rect 1055 1555 1095 1565
rect 1055 1285 1065 1555
rect 1085 1285 1095 1555
rect 1055 1275 1095 1285
rect 1155 1555 1195 1565
rect 1155 1285 1165 1555
rect 1185 1285 1195 1555
rect 1155 1275 1195 1285
rect 1255 1555 1295 1565
rect 1255 1285 1265 1555
rect 1285 1285 1295 1555
rect 1255 1275 1295 1285
rect 1355 1555 1395 1565
rect 1355 1285 1365 1555
rect 1385 1285 1395 1555
rect 1355 1275 1395 1285
rect 1455 1555 1495 1565
rect 1455 1285 1465 1555
rect 1485 1285 1495 1555
rect 1455 1275 1495 1285
rect 1555 1555 1595 1565
rect 1555 1285 1565 1555
rect 1585 1285 1595 1555
rect 1555 1275 1595 1285
rect 1655 1555 1695 1565
rect 1655 1285 1665 1555
rect 1685 1285 1695 1555
rect 1655 1275 1695 1285
rect 1755 1555 2085 1565
rect 1755 1285 1765 1555
rect 1785 1285 1815 1555
rect 2075 1285 2085 1555
rect 1755 1275 2085 1285
rect -45 1255 -5 1275
rect 165 1255 185 1275
rect 365 1255 385 1275
rect 765 1255 785 1275
rect 965 1255 985 1275
rect 1365 1255 1385 1275
rect 1565 1255 1585 1275
rect 1755 1255 1795 1275
rect -45 1245 50 1255
rect -45 1225 15 1245
rect 35 1225 50 1245
rect -45 1215 50 1225
rect 100 1245 1650 1255
rect 100 1225 115 1245
rect 135 1225 215 1245
rect 235 1225 315 1245
rect 335 1225 415 1245
rect 435 1225 515 1245
rect 535 1225 615 1245
rect 635 1225 715 1245
rect 735 1225 815 1245
rect 835 1225 915 1245
rect 935 1225 1015 1245
rect 1035 1225 1115 1245
rect 1135 1225 1215 1245
rect 1235 1225 1315 1245
rect 1335 1225 1415 1245
rect 1435 1225 1515 1245
rect 1535 1225 1615 1245
rect 1635 1225 1650 1245
rect 100 1215 1650 1225
rect 1700 1245 1795 1255
rect 1700 1225 1715 1245
rect 1735 1225 1795 1245
rect 1700 1215 1795 1225
rect 415 1175 1435 1195
rect -335 1165 -240 1175
rect -335 1145 -275 1165
rect -255 1145 -240 1165
rect -335 1135 -240 1145
rect -215 1165 390 1175
rect -215 1145 -175 1165
rect -155 1145 -75 1165
rect -55 1145 25 1165
rect 45 1145 125 1165
rect 145 1145 355 1165
rect 375 1145 390 1165
rect -215 1135 390 1145
rect -335 1105 -295 1135
rect -215 1115 -195 1135
rect -25 1115 -5 1135
rect 175 1115 195 1135
rect 415 1115 435 1175
rect 495 1135 1055 1155
rect 495 1115 515 1135
rect 1035 1115 1055 1135
rect 1415 1115 1435 1175
rect 1590 1165 1940 1175
rect 1590 1145 1605 1165
rect 1625 1145 1705 1165
rect 1725 1145 1805 1165
rect 1825 1145 1905 1165
rect 1925 1145 1940 1165
rect 1590 1135 1940 1145
rect 1990 1165 2085 1175
rect 1990 1145 2005 1165
rect 2025 1145 2085 1165
rect 1990 1135 2085 1145
rect 1655 1115 1675 1135
rect 1855 1115 1875 1135
rect -335 835 -325 1105
rect -305 835 -295 1105
rect -335 825 -295 835
rect -235 1105 -195 1115
rect -235 835 -225 1105
rect -205 835 -195 1105
rect -235 825 -195 835
rect -135 1105 -95 1115
rect -135 835 -125 1105
rect -105 835 -95 1105
rect -135 825 -95 835
rect -35 1105 5 1115
rect -35 835 -25 1105
rect -5 835 5 1105
rect -35 825 5 835
rect 65 1105 105 1115
rect 65 835 75 1105
rect 95 835 105 1105
rect 65 825 105 835
rect 165 1105 205 1115
rect 165 835 175 1105
rect 195 835 205 1105
rect 165 825 205 835
rect 245 1105 335 1115
rect 245 835 255 1105
rect 275 835 305 1105
rect 325 835 335 1105
rect 245 825 335 835
rect 395 1105 435 1115
rect 395 835 405 1105
rect 425 835 435 1105
rect 395 825 435 835
rect 475 1105 515 1115
rect 475 835 485 1105
rect 505 835 515 1105
rect 475 825 515 835
rect 575 1105 615 1115
rect 575 835 585 1105
rect 605 835 615 1105
rect 575 825 615 835
rect 675 1105 715 1115
rect 675 835 685 1105
rect 705 835 715 1105
rect 675 825 715 835
rect 755 1105 795 1115
rect 755 835 765 1105
rect 785 835 795 1105
rect 755 825 795 835
rect 855 1105 895 1115
rect 855 835 865 1105
rect 885 835 895 1105
rect 855 825 895 835
rect 955 1105 995 1115
rect 955 835 965 1105
rect 985 835 995 1105
rect 955 825 995 835
rect 1035 1105 1075 1115
rect 1035 835 1045 1105
rect 1065 835 1075 1105
rect 1035 825 1075 835
rect 1135 1105 1175 1115
rect 1135 835 1145 1105
rect 1165 835 1175 1105
rect 1135 825 1175 835
rect 1235 1105 1275 1115
rect 1235 835 1245 1105
rect 1265 835 1275 1105
rect 1235 825 1275 835
rect 1315 1105 1355 1115
rect 1315 835 1325 1105
rect 1345 835 1355 1105
rect 1315 825 1355 835
rect 1415 1105 1505 1115
rect 1415 835 1425 1105
rect 1445 835 1475 1105
rect 1495 835 1505 1105
rect 1415 825 1505 835
rect 1545 1105 1585 1115
rect 1545 835 1555 1105
rect 1575 835 1585 1105
rect 1545 825 1585 835
rect 1645 1105 1685 1115
rect 1645 835 1655 1105
rect 1675 835 1685 1105
rect 1645 825 1685 835
rect 1745 1105 1785 1115
rect 1745 835 1755 1105
rect 1775 835 1785 1105
rect 1745 825 1785 835
rect 1845 1105 1885 1115
rect 1845 835 1855 1105
rect 1875 835 1885 1105
rect 1845 825 1885 835
rect 1945 1105 1985 1115
rect 1945 835 1955 1105
rect 1975 835 1985 1105
rect 1945 825 1985 835
rect 2045 1105 2085 1135
rect 2045 835 2055 1105
rect 2075 835 2085 1105
rect 2045 825 2085 835
rect 695 785 715 825
rect 765 805 785 825
rect 965 805 985 825
rect 1315 805 1335 825
rect 765 785 1335 805
rect 1555 805 1575 825
rect 1755 805 1775 825
rect 1955 805 1975 825
rect 1555 785 1975 805
rect 695 725 715 765
rect 765 745 1335 765
rect 765 725 785 745
rect 965 725 985 745
rect 1315 725 1335 745
rect 1555 745 1975 765
rect 1555 725 1575 745
rect 1755 725 1775 745
rect 1955 725 1975 745
rect -335 715 -295 725
rect -335 445 -325 715
rect -305 445 -295 715
rect -335 415 -295 445
rect -235 715 -195 725
rect -235 445 -225 715
rect -205 445 -195 715
rect -235 435 -195 445
rect -135 715 -95 725
rect -135 445 -125 715
rect -105 445 -95 715
rect -135 435 -95 445
rect -35 715 5 725
rect -35 445 -25 715
rect -5 445 5 715
rect -35 435 5 445
rect 65 715 105 725
rect 65 445 75 715
rect 95 445 105 715
rect 65 435 105 445
rect 165 715 205 725
rect 165 445 175 715
rect 195 445 205 715
rect 165 435 205 445
rect 245 715 335 725
rect 245 445 255 715
rect 275 445 305 715
rect 325 445 335 715
rect 245 435 335 445
rect 395 715 435 725
rect 395 445 405 715
rect 425 445 435 715
rect 395 435 435 445
rect 475 715 515 725
rect 475 445 485 715
rect 505 445 515 715
rect 475 435 515 445
rect 575 715 615 725
rect 575 445 585 715
rect 605 445 615 715
rect 575 435 615 445
rect 675 715 715 725
rect 675 445 685 715
rect 705 445 715 715
rect 675 435 715 445
rect 755 715 795 725
rect 755 445 765 715
rect 785 445 795 715
rect 755 435 795 445
rect 855 715 895 725
rect 855 445 865 715
rect 885 445 895 715
rect 855 435 895 445
rect 955 715 995 725
rect 955 445 965 715
rect 985 445 995 715
rect 955 435 995 445
rect 1035 715 1075 725
rect 1035 445 1045 715
rect 1065 445 1075 715
rect 1035 435 1075 445
rect 1135 715 1175 725
rect 1135 445 1145 715
rect 1165 445 1175 715
rect 1135 435 1175 445
rect 1235 715 1275 725
rect 1235 445 1245 715
rect 1265 445 1275 715
rect 1235 435 1275 445
rect 1315 715 1355 725
rect 1315 445 1325 715
rect 1345 445 1355 715
rect 1315 435 1355 445
rect 1415 715 1505 725
rect 1415 445 1425 715
rect 1445 445 1475 715
rect 1495 445 1505 715
rect 1415 435 1505 445
rect 1545 715 1585 725
rect 1545 445 1555 715
rect 1575 445 1585 715
rect 1545 435 1585 445
rect 1645 715 1685 725
rect 1645 445 1655 715
rect 1675 445 1685 715
rect 1645 435 1685 445
rect 1745 715 1785 725
rect 1745 445 1755 715
rect 1775 445 1785 715
rect 1745 435 1785 445
rect 1845 715 1885 725
rect 1845 445 1855 715
rect 1875 445 1885 715
rect 1845 435 1885 445
rect 1945 715 1985 725
rect 1945 445 1955 715
rect 1975 445 1985 715
rect 1945 435 1985 445
rect 2045 715 2085 725
rect 2045 445 2055 715
rect 2075 445 2085 715
rect -215 415 -195 435
rect -25 415 -5 435
rect 175 415 195 435
rect -335 405 -240 415
rect -335 385 -275 405
rect -255 385 -240 405
rect -335 375 -240 385
rect -215 405 390 415
rect -215 385 -175 405
rect -155 385 -75 405
rect -55 385 25 405
rect 45 385 125 405
rect 145 385 355 405
rect 375 385 390 405
rect -215 375 390 385
rect 415 375 435 435
rect 495 415 515 435
rect 1035 415 1055 435
rect 495 395 1055 415
rect 1415 375 1435 435
rect 1655 415 1675 435
rect 1855 415 1875 435
rect 2045 415 2085 445
rect 1590 405 1940 415
rect 1590 385 1605 405
rect 1625 385 1705 405
rect 1725 385 1805 405
rect 1825 385 1905 405
rect 1925 385 1940 405
rect 1590 375 1940 385
rect 1990 405 2085 415
rect 1990 385 2005 405
rect 2025 385 2085 405
rect 1990 375 2085 385
rect 415 355 1435 375
rect -45 325 50 335
rect -45 305 15 325
rect 35 305 50 325
rect -45 295 50 305
rect 100 325 1650 335
rect 100 305 115 325
rect 135 305 215 325
rect 235 305 315 325
rect 335 305 415 325
rect 435 305 515 325
rect 535 305 615 325
rect 635 305 715 325
rect 735 305 815 325
rect 835 305 915 325
rect 935 305 1015 325
rect 1035 305 1115 325
rect 1135 305 1215 325
rect 1235 305 1315 325
rect 1335 305 1415 325
rect 1435 305 1515 325
rect 1535 305 1615 325
rect 1635 305 1650 325
rect 100 295 1650 305
rect 1700 325 1795 335
rect 1700 305 1715 325
rect 1735 305 1795 325
rect 1700 295 1795 305
rect -45 275 -5 295
rect 165 275 185 295
rect 365 275 385 295
rect 765 275 785 295
rect 965 275 985 295
rect 1365 275 1385 295
rect 1565 275 1585 295
rect 1755 275 1795 295
rect -335 265 -5 275
rect -335 -5 -325 265
rect -65 -5 -35 265
rect -15 -5 -5 265
rect -335 -15 -5 -5
rect 55 265 95 275
rect 55 -5 65 265
rect 85 -5 95 265
rect 55 -15 95 -5
rect 155 265 195 275
rect 155 -5 165 265
rect 185 -5 195 265
rect 155 -15 195 -5
rect 255 265 295 275
rect 255 -5 265 265
rect 285 -5 295 265
rect 255 -15 295 -5
rect 355 265 395 275
rect 355 -5 365 265
rect 385 -5 395 265
rect 355 -15 395 -5
rect 455 265 495 275
rect 455 -5 465 265
rect 485 -5 495 265
rect 455 -15 495 -5
rect 555 265 595 275
rect 555 -5 565 265
rect 585 -5 595 265
rect 555 -15 595 -5
rect 655 265 695 275
rect 655 -5 665 265
rect 685 -5 695 265
rect 655 -15 695 -5
rect 755 265 795 275
rect 755 -5 765 265
rect 785 -5 795 265
rect 755 -15 795 -5
rect 855 265 895 275
rect 855 -5 865 265
rect 885 -5 895 265
rect 855 -15 895 -5
rect 955 265 995 275
rect 955 -5 965 265
rect 985 -5 995 265
rect 955 -15 995 -5
rect 1055 265 1095 275
rect 1055 -5 1065 265
rect 1085 -5 1095 265
rect 1055 -15 1095 -5
rect 1155 265 1195 275
rect 1155 -5 1165 265
rect 1185 -5 1195 265
rect 1155 -15 1195 -5
rect 1255 265 1295 275
rect 1255 -5 1265 265
rect 1285 -5 1295 265
rect 1255 -15 1295 -5
rect 1355 265 1395 275
rect 1355 -5 1365 265
rect 1385 -5 1395 265
rect 1355 -15 1395 -5
rect 1455 265 1495 275
rect 1455 -5 1465 265
rect 1485 -5 1495 265
rect 1455 -15 1495 -5
rect 1555 265 1595 275
rect 1555 -5 1565 265
rect 1585 -5 1595 265
rect 1555 -15 1595 -5
rect 1655 265 1695 275
rect 1655 -5 1665 265
rect 1685 -5 1695 265
rect 1655 -15 1695 -5
rect 1755 265 2085 275
rect 1755 -5 1765 265
rect 1785 -5 1815 265
rect 2075 -5 2085 265
rect 1755 -15 2085 -5
rect 65 -35 85 -15
rect 265 -35 285 -15
rect 465 -35 485 -15
rect 665 -35 685 -15
rect 865 -35 885 -15
rect 1065 -35 1085 -15
rect 1265 -35 1285 -15
rect 1465 -35 1485 -15
rect 1665 -35 1685 -15
rect 65 -55 1685 -35
<< viali >>
rect -325 1285 -65 1555
rect -35 1285 -15 1555
rect 565 1285 585 1555
rect 1165 1285 1185 1555
rect 1765 1285 1785 1555
rect 1815 1285 2075 1555
rect -325 835 -305 1105
rect -125 835 -105 1105
rect 75 835 95 1105
rect 255 835 275 1105
rect 305 835 325 1105
rect 865 835 885 1105
rect 1245 835 1265 1105
rect 1425 835 1445 1105
rect 1475 835 1495 1105
rect 2055 835 2075 1105
rect -325 445 -305 715
rect -125 445 -105 715
rect 75 445 95 715
rect 255 445 275 715
rect 305 445 325 715
rect 865 445 885 715
rect 1245 445 1265 715
rect 1425 445 1445 715
rect 1475 445 1495 715
rect 2055 445 2075 715
rect -325 -5 -65 265
rect -35 -5 -15 265
rect 565 -5 585 265
rect 1165 -5 1185 265
rect 1765 -5 1785 265
rect 1815 -5 2075 265
<< metal1 >>
rect -45 1555 -5 1565
rect -45 1285 -35 1555
rect -15 1285 -5 1555
rect -45 1275 -5 1285
rect 555 1555 595 1565
rect 555 1285 565 1555
rect 585 1285 595 1555
rect 555 1275 595 1285
rect 1155 1555 1195 1565
rect 1155 1285 1165 1555
rect 1185 1285 1195 1555
rect 1155 1275 1195 1285
rect 1755 1555 1795 1565
rect 1755 1285 1765 1555
rect 1785 1285 1795 1555
rect 1755 1275 1795 1285
rect -335 1105 -295 1115
rect 2045 1105 2085 1115
rect -335 835 -325 1105
rect -305 835 -295 1105
rect 2045 835 2055 1105
rect 2075 835 2085 1105
rect -335 825 -295 835
rect 2045 825 2085 835
rect -335 715 -295 725
rect 2045 715 2085 725
rect -335 445 -325 715
rect -305 445 -295 715
rect 2045 445 2055 715
rect 2075 445 2085 715
rect -335 435 -295 445
rect 2045 435 2085 445
rect -45 265 -5 275
rect -45 -5 -35 265
rect -15 -5 -5 265
rect -45 -15 -5 -5
rect 555 265 595 275
rect 555 -5 565 265
rect 585 -5 595 265
rect 555 -15 595 -5
rect 1155 265 1195 275
rect 1155 -5 1165 265
rect 1185 -5 1195 265
rect 1155 -15 1195 -5
rect 1755 265 1795 275
rect 1755 -5 1765 265
rect 1785 -5 1795 265
rect 1755 -15 1795 -5
<< end >>
