magic
tech sky130A
timestamp 1697129809
<< nmos >>
rect 0 -20 50 280
rect 100 -20 150 280
rect 200 -20 250 280
rect 300 -20 350 280
rect 400 -20 450 280
rect 500 -20 550 280
rect 600 -20 650 280
rect 700 -20 750 280
rect 800 -20 850 280
rect 900 -20 950 280
rect 1000 -20 1050 280
rect 1100 -20 1150 280
rect 1200 -20 1250 280
rect 1300 -20 1350 280
rect 1400 -20 1450 280
rect 1500 -20 1550 280
rect 1600 -20 1650 280
rect 1700 -20 1750 280
<< ndiff >>
rect -50 265 0 280
rect -50 -5 -35 265
rect -15 -5 0 265
rect -50 -20 0 -5
rect 50 265 100 280
rect 50 -5 65 265
rect 85 -5 100 265
rect 50 -20 100 -5
rect 150 265 200 280
rect 150 -5 165 265
rect 185 -5 200 265
rect 150 -20 200 -5
rect 250 265 300 280
rect 250 -5 265 265
rect 285 -5 300 265
rect 250 -20 300 -5
rect 350 265 400 280
rect 350 -5 365 265
rect 385 -5 400 265
rect 350 -20 400 -5
rect 450 265 500 280
rect 450 -5 465 265
rect 485 -5 500 265
rect 450 -20 500 -5
rect 550 265 600 280
rect 550 -5 565 265
rect 585 -5 600 265
rect 550 -20 600 -5
rect 650 265 700 280
rect 650 -5 665 265
rect 685 -5 700 265
rect 650 -20 700 -5
rect 750 265 800 280
rect 750 -5 765 265
rect 785 -5 800 265
rect 750 -20 800 -5
rect 850 265 900 280
rect 850 -5 865 265
rect 885 -5 900 265
rect 850 -20 900 -5
rect 950 265 1000 280
rect 950 -5 965 265
rect 985 -5 1000 265
rect 950 -20 1000 -5
rect 1050 265 1100 280
rect 1050 -5 1065 265
rect 1085 -5 1100 265
rect 1050 -20 1100 -5
rect 1150 265 1200 280
rect 1150 -5 1165 265
rect 1185 -5 1200 265
rect 1150 -20 1200 -5
rect 1250 265 1300 280
rect 1250 -5 1265 265
rect 1285 -5 1300 265
rect 1250 -20 1300 -5
rect 1350 265 1400 280
rect 1350 -5 1365 265
rect 1385 -5 1400 265
rect 1350 -20 1400 -5
rect 1450 265 1500 280
rect 1450 -5 1465 265
rect 1485 -5 1500 265
rect 1450 -20 1500 -5
rect 1550 265 1600 280
rect 1550 -5 1565 265
rect 1585 -5 1600 265
rect 1550 -20 1600 -5
rect 1650 265 1700 280
rect 1650 -5 1665 265
rect 1685 -5 1700 265
rect 1650 -20 1700 -5
rect 1750 265 1800 280
rect 1750 -5 1765 265
rect 1785 -5 1800 265
rect 1750 -20 1800 -5
<< ndiffc >>
rect -35 -5 -15 265
rect 65 -5 85 265
rect 165 -5 185 265
rect 265 -5 285 265
rect 365 -5 385 265
rect 465 -5 485 265
rect 565 -5 585 265
rect 665 -5 685 265
rect 765 -5 785 265
rect 865 -5 885 265
rect 965 -5 985 265
rect 1065 -5 1085 265
rect 1165 -5 1185 265
rect 1265 -5 1285 265
rect 1365 -5 1385 265
rect 1465 -5 1485 265
rect 1565 -5 1585 265
rect 1665 -5 1685 265
rect 1765 -5 1785 265
<< poly >>
rect 0 325 50 335
rect 0 305 15 325
rect 35 305 50 325
rect 0 280 50 305
rect 100 325 150 335
rect 100 305 115 325
rect 135 305 150 325
rect 100 280 150 305
rect 200 325 250 335
rect 200 305 215 325
rect 235 305 250 325
rect 200 280 250 305
rect 300 325 350 335
rect 300 305 315 325
rect 335 305 350 325
rect 300 280 350 305
rect 400 325 450 335
rect 400 305 415 325
rect 435 305 450 325
rect 400 280 450 305
rect 500 325 550 335
rect 500 305 515 325
rect 535 305 550 325
rect 500 280 550 305
rect 600 325 650 335
rect 600 305 615 325
rect 635 305 650 325
rect 600 280 650 305
rect 700 325 750 335
rect 700 305 715 325
rect 735 305 750 325
rect 700 280 750 305
rect 800 325 850 335
rect 800 305 815 325
rect 835 305 850 325
rect 800 280 850 305
rect 900 325 950 335
rect 900 305 915 325
rect 935 305 950 325
rect 900 280 950 305
rect 1000 325 1050 335
rect 1000 305 1015 325
rect 1035 305 1050 325
rect 1000 280 1050 305
rect 1100 325 1150 335
rect 1100 305 1115 325
rect 1135 305 1150 325
rect 1100 280 1150 305
rect 1200 325 1250 335
rect 1200 305 1215 325
rect 1235 305 1250 325
rect 1200 280 1250 305
rect 1300 325 1350 335
rect 1300 305 1315 325
rect 1335 305 1350 325
rect 1300 280 1350 305
rect 1400 325 1450 335
rect 1400 305 1415 325
rect 1435 305 1450 325
rect 1400 280 1450 305
rect 1500 325 1550 335
rect 1500 305 1515 325
rect 1535 305 1550 325
rect 1500 280 1550 305
rect 1600 325 1650 335
rect 1600 305 1615 325
rect 1635 305 1650 325
rect 1600 280 1650 305
rect 1700 325 1750 335
rect 1700 305 1715 325
rect 1735 305 1750 325
rect 1700 280 1750 305
rect 0 -35 50 -20
rect 100 -35 150 -20
rect 200 -35 250 -20
rect 300 -35 350 -20
rect 400 -35 450 -20
rect 500 -35 550 -20
rect 600 -35 650 -20
rect 700 -35 750 -20
rect 800 -35 850 -20
rect 900 -35 950 -20
rect 1000 -35 1050 -20
rect 1100 -35 1150 -20
rect 1200 -35 1250 -20
rect 1300 -35 1350 -20
rect 1400 -35 1450 -20
rect 1500 -35 1550 -20
rect 1600 -35 1650 -20
rect 1700 -35 1750 -20
<< polycont >>
rect 15 305 35 325
rect 115 305 135 325
rect 215 305 235 325
rect 315 305 335 325
rect 415 305 435 325
rect 515 305 535 325
rect 615 305 635 325
rect 715 305 735 325
rect 815 305 835 325
rect 915 305 935 325
rect 1015 305 1035 325
rect 1115 305 1135 325
rect 1215 305 1235 325
rect 1315 305 1335 325
rect 1415 305 1435 325
rect 1515 305 1535 325
rect 1615 305 1635 325
rect 1715 305 1735 325
<< locali >>
rect -45 325 50 335
rect -45 305 15 325
rect 35 305 50 325
rect -45 295 50 305
rect 100 325 1650 335
rect 100 305 115 325
rect 135 305 215 325
rect 235 305 315 325
rect 335 305 415 325
rect 435 305 515 325
rect 535 305 615 325
rect 635 305 715 325
rect 735 305 815 325
rect 835 305 915 325
rect 935 305 1015 325
rect 1035 305 1115 325
rect 1135 305 1215 325
rect 1235 305 1315 325
rect 1335 305 1415 325
rect 1435 305 1515 325
rect 1535 305 1615 325
rect 1635 305 1650 325
rect 100 295 1650 305
rect 1700 325 1795 335
rect 1700 305 1715 325
rect 1735 305 1795 325
rect 1700 295 1795 305
rect -45 265 -5 295
rect 165 275 185 295
rect 365 275 385 295
rect 765 275 785 295
rect 965 275 985 295
rect 1365 275 1385 295
rect 1565 275 1585 295
rect -45 -5 -35 265
rect -15 -5 -5 265
rect -45 -15 -5 -5
rect 55 265 95 275
rect 55 -5 65 265
rect 85 -5 95 265
rect 55 -15 95 -5
rect 155 265 195 275
rect 155 -5 165 265
rect 185 -5 195 265
rect 155 -15 195 -5
rect 255 265 295 275
rect 255 -5 265 265
rect 285 -5 295 265
rect 255 -15 295 -5
rect 355 265 395 275
rect 355 -5 365 265
rect 385 -5 395 265
rect 355 -15 395 -5
rect 455 265 495 275
rect 455 -5 465 265
rect 485 -5 495 265
rect 455 -15 495 -5
rect 555 265 595 275
rect 555 -5 565 265
rect 585 -5 595 265
rect 555 -15 595 -5
rect 655 265 695 275
rect 655 -5 665 265
rect 685 -5 695 265
rect 655 -15 695 -5
rect 755 265 795 275
rect 755 -5 765 265
rect 785 -5 795 265
rect 755 -15 795 -5
rect 855 265 895 275
rect 855 -5 865 265
rect 885 -5 895 265
rect 855 -15 895 -5
rect 955 265 995 275
rect 955 -5 965 265
rect 985 -5 995 265
rect 955 -15 995 -5
rect 1055 265 1095 275
rect 1055 -5 1065 265
rect 1085 -5 1095 265
rect 1055 -15 1095 -5
rect 1155 265 1195 275
rect 1155 -5 1165 265
rect 1185 -5 1195 265
rect 1155 -15 1195 -5
rect 1255 265 1295 275
rect 1255 -5 1265 265
rect 1285 -5 1295 265
rect 1255 -15 1295 -5
rect 1355 265 1395 275
rect 1355 -5 1365 265
rect 1385 -5 1395 265
rect 1355 -15 1395 -5
rect 1455 265 1495 275
rect 1455 -5 1465 265
rect 1485 -5 1495 265
rect 1455 -15 1495 -5
rect 1555 265 1595 275
rect 1555 -5 1565 265
rect 1585 -5 1595 265
rect 1555 -15 1595 -5
rect 1655 265 1695 275
rect 1655 -5 1665 265
rect 1685 -5 1695 265
rect 1655 -15 1695 -5
rect 1755 265 1795 295
rect 1755 -5 1765 265
rect 1785 -5 1795 265
rect 1755 -15 1795 -5
rect 65 -35 85 -15
rect 265 -35 285 -15
rect 465 -35 485 -15
rect 665 -35 685 -15
rect 865 -35 885 -15
rect 1065 -35 1085 -15
rect 1265 -35 1285 -15
rect 1465 -35 1485 -15
rect 1665 -35 1685 -15
rect 65 -55 1685 -35
<< viali >>
rect -35 -5 -15 265
rect 565 -5 585 265
rect 1165 -5 1185 265
rect 1765 -5 1785 265
<< metal1 >>
rect -45 265 -5 275
rect -45 -5 -35 265
rect -15 -5 -5 265
rect -45 -15 -5 -5
rect 555 265 595 275
rect 555 -5 565 265
rect 585 -5 595 265
rect 555 -15 595 -5
rect 1155 265 1195 275
rect 1155 -5 1165 265
rect 1185 -5 1195 265
rect 1155 -15 1195 -5
rect 1755 265 1795 275
rect 1755 -5 1765 265
rect 1785 -5 1795 265
rect 1755 -15 1795 -5
<< end >>
