magic
tech sky130A
timestamp 1693857689
<< nwell >>
rect -120 135 200 275
<< nmos >>
rect 0 0 15 100
rect 65 0 80 100
<< pmos >>
rect 0 155 15 255
rect 65 155 80 255
<< ndiff >>
rect -55 85 0 100
rect -55 15 -35 85
rect -15 15 0 85
rect -55 0 0 15
rect 15 0 65 100
rect 80 85 130 100
rect 80 15 95 85
rect 115 15 130 85
rect 80 0 130 15
<< pdiff >>
rect -50 240 0 255
rect -50 170 -35 240
rect -15 170 0 240
rect -50 155 0 170
rect 15 240 65 255
rect 15 170 30 240
rect 50 170 65 240
rect 15 155 65 170
rect 80 240 130 255
rect 80 170 95 240
rect 115 170 130 240
rect 80 155 130 170
<< ndiffc >>
rect -35 15 -15 85
rect 95 15 115 85
<< pdiffc >>
rect -35 170 -15 240
rect 30 170 50 240
rect 95 170 115 240
<< psubdiff >>
rect -110 85 -55 100
rect -110 15 -95 85
rect -75 15 -55 85
rect -110 0 -55 15
rect 130 85 180 100
rect 130 15 145 85
rect 165 15 180 85
rect 130 0 180 15
<< nsubdiff >>
rect -100 240 -50 255
rect -100 170 -85 240
rect -65 170 -50 240
rect -100 155 -50 170
rect 130 240 180 255
rect 130 170 145 240
rect 165 170 180 240
rect 130 155 180 170
<< psubdiffcont >>
rect -95 15 -75 85
rect 145 15 165 85
<< nsubdiffcont >>
rect -85 170 -65 240
rect 145 170 165 240
<< poly >>
rect 0 255 15 270
rect 65 255 80 270
rect 0 100 15 155
rect 65 100 80 155
rect 0 -15 15 0
rect -40 -25 15 -15
rect -40 -45 -30 -25
rect -10 -35 15 -25
rect -10 -45 0 -35
rect -40 -55 0 -45
rect 65 -55 80 0
rect 40 -65 80 -55
rect 40 -85 50 -65
rect 70 -85 80 -65
rect 40 -95 80 -85
<< polycont >>
rect -30 -45 -10 -25
rect 50 -85 70 -65
<< locali >>
rect -95 240 -5 250
rect -95 170 -85 240
rect -65 170 -35 240
rect -15 170 -5 240
rect -95 160 -5 170
rect 20 240 60 250
rect 20 170 30 240
rect 50 170 60 240
rect 20 160 60 170
rect 85 240 175 250
rect 85 170 95 240
rect 115 170 145 240
rect 165 170 175 240
rect 85 160 175 170
rect 20 95 40 160
rect -105 85 -65 95
rect -105 15 -95 85
rect -75 15 -65 85
rect -105 5 -65 15
rect -45 85 40 95
rect -45 15 -35 85
rect -15 75 40 85
rect -15 15 -5 75
rect -45 5 -5 15
rect 20 -15 40 75
rect 85 85 175 95
rect 85 15 95 85
rect 115 15 145 85
rect 165 15 175 85
rect 85 5 175 15
rect -120 -25 0 -15
rect -120 -35 -30 -25
rect -40 -45 -30 -35
rect -10 -45 0 -25
rect 20 -35 200 -15
rect -40 -55 0 -45
rect 40 -65 80 -55
rect 40 -75 50 -65
rect -120 -85 50 -75
rect 70 -85 80 -65
rect -120 -95 80 -85
<< viali >>
rect -85 170 -65 240
rect -35 170 -15 240
rect 95 170 115 240
rect 145 170 165 240
rect -95 15 -75 85
rect 95 15 115 85
rect 145 15 165 85
<< metal1 >>
rect -120 240 200 255
rect -120 170 -85 240
rect -65 170 -35 240
rect -15 170 95 240
rect 115 170 145 240
rect 165 170 200 240
rect -120 155 200 170
rect -120 85 200 100
rect -120 15 -95 85
rect -75 15 95 85
rect 115 15 145 85
rect 165 15 200 85
rect -120 0 200 15
<< labels >>
rlabel locali -120 -25 -120 -25 7 A
port 1 w
rlabel locali -120 -85 -120 -85 7 B
port 2 w
rlabel metal1 -120 205 -120 205 7 VP
port 4 w
rlabel metal1 -120 50 -120 50 7 VN
port 5 w
rlabel locali 200 -25 200 -25 3 Y
port 3 e
<< end >>
