magic
tech sky130A
timestamp 1697158498
<< nwell >>
rect -360 1175 2110 1590
rect -760 800 2110 1175
<< nmos >>
rect -290 410 -240 710
rect -190 410 -140 710
rect -90 410 -40 710
rect 10 410 60 710
rect 110 410 160 710
rect 340 410 390 710
rect 520 410 570 710
rect 620 410 670 710
rect 800 410 850 710
rect 900 410 950 710
rect 1080 410 1130 710
rect 1180 410 1230 710
rect 1360 410 1410 710
rect 1590 395 1640 695
rect 1690 395 1740 695
rect 1790 395 1840 695
rect 1890 395 1940 695
rect 1990 395 2040 695
rect 0 -40 50 260
rect 100 -40 150 260
rect 200 -40 250 260
rect 300 -40 350 260
rect 400 -40 450 260
rect 500 -40 550 260
rect 600 -40 650 260
rect 700 -40 750 260
rect 800 -40 850 260
rect 900 -40 950 260
rect 1000 -40 1050 260
rect 1100 -40 1150 260
rect 1200 -40 1250 260
rect 1300 -40 1350 260
rect 1400 -40 1450 260
rect 1500 -40 1550 260
rect 1600 -40 1650 260
rect 1700 -40 1750 260
<< pmos >>
rect 0 1270 50 1570
rect 100 1270 150 1570
rect 200 1270 250 1570
rect 300 1270 350 1570
rect 400 1270 450 1570
rect 500 1270 550 1570
rect 600 1270 650 1570
rect 700 1270 750 1570
rect 800 1270 850 1570
rect 900 1270 950 1570
rect 1000 1270 1050 1570
rect 1100 1270 1150 1570
rect 1200 1270 1250 1570
rect 1300 1270 1350 1570
rect 1400 1270 1450 1570
rect 1500 1270 1550 1570
rect 1600 1270 1650 1570
rect 1700 1270 1750 1570
rect -690 820 -640 1120
rect -590 820 -540 1120
rect -490 820 -440 1120
rect -390 820 -340 1120
rect -290 820 -240 1120
rect -190 820 -140 1120
rect -90 820 -40 1120
rect 10 820 60 1120
rect 110 820 160 1120
rect 340 820 390 1120
rect 520 820 570 1120
rect 620 820 670 1120
rect 800 820 850 1120
rect 900 820 950 1120
rect 1080 820 1130 1120
rect 1180 820 1230 1120
rect 1360 820 1410 1120
rect 1590 835 1640 1135
rect 1690 835 1740 1135
rect 1790 835 1840 1135
rect 1890 835 1940 1135
rect 1990 835 2040 1135
<< ndiff >>
rect -340 695 -290 710
rect -340 425 -325 695
rect -305 425 -290 695
rect -340 410 -290 425
rect -240 695 -190 710
rect -240 425 -225 695
rect -205 425 -190 695
rect -240 410 -190 425
rect -140 695 -90 710
rect -140 425 -125 695
rect -105 425 -90 695
rect -140 410 -90 425
rect -40 695 10 710
rect -40 425 -25 695
rect -5 425 10 695
rect -40 410 10 425
rect 60 695 110 710
rect 60 425 75 695
rect 95 425 110 695
rect 60 410 110 425
rect 160 695 210 710
rect 160 425 175 695
rect 195 425 210 695
rect 160 410 210 425
rect 290 695 340 710
rect 290 425 305 695
rect 325 425 340 695
rect 290 410 340 425
rect 390 695 440 710
rect 390 425 405 695
rect 425 425 440 695
rect 390 410 440 425
rect 470 695 520 710
rect 470 425 485 695
rect 505 425 520 695
rect 470 410 520 425
rect 570 695 620 710
rect 570 425 585 695
rect 605 425 620 695
rect 570 410 620 425
rect 670 695 720 710
rect 670 425 685 695
rect 705 425 720 695
rect 670 410 720 425
rect 750 695 800 710
rect 750 425 765 695
rect 785 425 800 695
rect 750 410 800 425
rect 850 695 900 710
rect 850 425 865 695
rect 885 425 900 695
rect 850 410 900 425
rect 950 695 1000 710
rect 950 425 965 695
rect 985 425 1000 695
rect 950 410 1000 425
rect 1030 695 1080 710
rect 1030 425 1045 695
rect 1065 425 1080 695
rect 1030 410 1080 425
rect 1130 695 1180 710
rect 1130 425 1145 695
rect 1165 425 1180 695
rect 1130 410 1180 425
rect 1230 695 1280 710
rect 1230 425 1245 695
rect 1265 425 1280 695
rect 1230 410 1280 425
rect 1310 695 1360 710
rect 1310 425 1325 695
rect 1345 425 1360 695
rect 1310 410 1360 425
rect 1410 695 1460 710
rect 1410 425 1425 695
rect 1445 425 1460 695
rect 1410 410 1460 425
rect 1540 680 1590 695
rect 1540 410 1555 680
rect 1575 410 1590 680
rect 1540 395 1590 410
rect 1640 680 1690 695
rect 1640 410 1655 680
rect 1675 410 1690 680
rect 1640 395 1690 410
rect 1740 680 1790 695
rect 1740 410 1755 680
rect 1775 410 1790 680
rect 1740 395 1790 410
rect 1840 680 1890 695
rect 1840 410 1855 680
rect 1875 410 1890 680
rect 1840 395 1890 410
rect 1940 680 1990 695
rect 1940 410 1955 680
rect 1975 410 1990 680
rect 1940 395 1990 410
rect 2040 680 2090 695
rect 2040 410 2055 680
rect 2075 410 2090 680
rect 2040 395 2090 410
rect -50 245 0 260
rect -50 -25 -35 245
rect -15 -25 0 245
rect -50 -40 0 -25
rect 50 245 100 260
rect 50 -25 65 245
rect 85 -25 100 245
rect 50 -40 100 -25
rect 150 245 200 260
rect 150 -25 165 245
rect 185 -25 200 245
rect 150 -40 200 -25
rect 250 245 300 260
rect 250 -25 265 245
rect 285 -25 300 245
rect 250 -40 300 -25
rect 350 245 400 260
rect 350 -25 365 245
rect 385 -25 400 245
rect 350 -40 400 -25
rect 450 245 500 260
rect 450 -25 465 245
rect 485 -25 500 245
rect 450 -40 500 -25
rect 550 245 600 260
rect 550 -25 565 245
rect 585 -25 600 245
rect 550 -40 600 -25
rect 650 245 700 260
rect 650 -25 665 245
rect 685 -25 700 245
rect 650 -40 700 -25
rect 750 245 800 260
rect 750 -25 765 245
rect 785 -25 800 245
rect 750 -40 800 -25
rect 850 245 900 260
rect 850 -25 865 245
rect 885 -25 900 245
rect 850 -40 900 -25
rect 950 245 1000 260
rect 950 -25 965 245
rect 985 -25 1000 245
rect 950 -40 1000 -25
rect 1050 245 1100 260
rect 1050 -25 1065 245
rect 1085 -25 1100 245
rect 1050 -40 1100 -25
rect 1150 245 1200 260
rect 1150 -25 1165 245
rect 1185 -25 1200 245
rect 1150 -40 1200 -25
rect 1250 245 1300 260
rect 1250 -25 1265 245
rect 1285 -25 1300 245
rect 1250 -40 1300 -25
rect 1350 245 1400 260
rect 1350 -25 1365 245
rect 1385 -25 1400 245
rect 1350 -40 1400 -25
rect 1450 245 1500 260
rect 1450 -25 1465 245
rect 1485 -25 1500 245
rect 1450 -40 1500 -25
rect 1550 245 1600 260
rect 1550 -25 1565 245
rect 1585 -25 1600 245
rect 1550 -40 1600 -25
rect 1650 245 1700 260
rect 1650 -25 1665 245
rect 1685 -25 1700 245
rect 1650 -40 1700 -25
rect 1750 245 1800 260
rect 1750 -25 1765 245
rect 1785 -25 1800 245
rect 1750 -40 1800 -25
<< pdiff >>
rect -50 1555 0 1570
rect -50 1285 -35 1555
rect -15 1285 0 1555
rect -50 1270 0 1285
rect 50 1555 100 1570
rect 50 1285 65 1555
rect 85 1285 100 1555
rect 50 1270 100 1285
rect 150 1555 200 1570
rect 150 1285 165 1555
rect 185 1285 200 1555
rect 150 1270 200 1285
rect 250 1555 300 1570
rect 250 1285 265 1555
rect 285 1285 300 1555
rect 250 1270 300 1285
rect 350 1555 400 1570
rect 350 1285 365 1555
rect 385 1285 400 1555
rect 350 1270 400 1285
rect 450 1555 500 1570
rect 450 1285 465 1555
rect 485 1285 500 1555
rect 450 1270 500 1285
rect 550 1555 600 1570
rect 550 1285 565 1555
rect 585 1285 600 1555
rect 550 1270 600 1285
rect 650 1555 700 1570
rect 650 1285 665 1555
rect 685 1285 700 1555
rect 650 1270 700 1285
rect 750 1555 800 1570
rect 750 1285 765 1555
rect 785 1285 800 1555
rect 750 1270 800 1285
rect 850 1555 900 1570
rect 850 1285 865 1555
rect 885 1285 900 1555
rect 850 1270 900 1285
rect 950 1555 1000 1570
rect 950 1285 965 1555
rect 985 1285 1000 1555
rect 950 1270 1000 1285
rect 1050 1555 1100 1570
rect 1050 1285 1065 1555
rect 1085 1285 1100 1555
rect 1050 1270 1100 1285
rect 1150 1555 1200 1570
rect 1150 1285 1165 1555
rect 1185 1285 1200 1555
rect 1150 1270 1200 1285
rect 1250 1555 1300 1570
rect 1250 1285 1265 1555
rect 1285 1285 1300 1555
rect 1250 1270 1300 1285
rect 1350 1555 1400 1570
rect 1350 1285 1365 1555
rect 1385 1285 1400 1555
rect 1350 1270 1400 1285
rect 1450 1555 1500 1570
rect 1450 1285 1465 1555
rect 1485 1285 1500 1555
rect 1450 1270 1500 1285
rect 1550 1555 1600 1570
rect 1550 1285 1565 1555
rect 1585 1285 1600 1555
rect 1550 1270 1600 1285
rect 1650 1555 1700 1570
rect 1650 1285 1665 1555
rect 1685 1285 1700 1555
rect 1650 1270 1700 1285
rect 1750 1555 1800 1570
rect 1750 1285 1765 1555
rect 1785 1285 1800 1555
rect 1750 1270 1800 1285
rect 1540 1120 1590 1135
rect -740 1105 -690 1120
rect -740 835 -725 1105
rect -705 835 -690 1105
rect -740 820 -690 835
rect -640 1105 -590 1120
rect -640 835 -625 1105
rect -605 835 -590 1105
rect -640 820 -590 835
rect -540 1105 -490 1120
rect -540 835 -525 1105
rect -505 835 -490 1105
rect -540 820 -490 835
rect -440 1105 -390 1120
rect -440 835 -425 1105
rect -405 835 -390 1105
rect -440 820 -390 835
rect -340 1105 -290 1120
rect -340 835 -325 1105
rect -305 835 -290 1105
rect -340 820 -290 835
rect -240 1105 -190 1120
rect -240 835 -225 1105
rect -205 835 -190 1105
rect -240 820 -190 835
rect -140 1105 -90 1120
rect -140 835 -125 1105
rect -105 835 -90 1105
rect -140 820 -90 835
rect -40 1105 10 1120
rect -40 835 -25 1105
rect -5 835 10 1105
rect -40 820 10 835
rect 60 1105 110 1120
rect 60 835 75 1105
rect 95 835 110 1105
rect 60 820 110 835
rect 160 1105 210 1120
rect 160 835 175 1105
rect 195 835 210 1105
rect 160 820 210 835
rect 290 1105 340 1120
rect 290 835 305 1105
rect 325 835 340 1105
rect 290 820 340 835
rect 390 1105 440 1120
rect 390 835 405 1105
rect 425 835 440 1105
rect 390 820 440 835
rect 470 1105 520 1120
rect 470 835 485 1105
rect 505 835 520 1105
rect 470 820 520 835
rect 570 1105 620 1120
rect 570 835 585 1105
rect 605 835 620 1105
rect 570 820 620 835
rect 670 1105 720 1120
rect 670 835 685 1105
rect 705 835 720 1105
rect 670 820 720 835
rect 750 1105 800 1120
rect 750 835 765 1105
rect 785 835 800 1105
rect 750 820 800 835
rect 850 1105 900 1120
rect 850 835 865 1105
rect 885 835 900 1105
rect 850 820 900 835
rect 950 1105 1000 1120
rect 950 835 965 1105
rect 985 835 1000 1105
rect 950 820 1000 835
rect 1030 1105 1080 1120
rect 1030 835 1045 1105
rect 1065 835 1080 1105
rect 1030 820 1080 835
rect 1130 1105 1180 1120
rect 1130 835 1145 1105
rect 1165 835 1180 1105
rect 1130 820 1180 835
rect 1230 1105 1280 1120
rect 1230 835 1245 1105
rect 1265 835 1280 1105
rect 1230 820 1280 835
rect 1310 1105 1360 1120
rect 1310 835 1325 1105
rect 1345 835 1360 1105
rect 1310 820 1360 835
rect 1410 1105 1460 1120
rect 1410 835 1425 1105
rect 1445 835 1460 1105
rect 1540 850 1555 1120
rect 1575 850 1590 1120
rect 1540 835 1590 850
rect 1640 1120 1690 1135
rect 1640 850 1655 1120
rect 1675 850 1690 1120
rect 1640 835 1690 850
rect 1740 1120 1790 1135
rect 1740 850 1755 1120
rect 1775 850 1790 1120
rect 1740 835 1790 850
rect 1840 1120 1890 1135
rect 1840 850 1855 1120
rect 1875 850 1890 1120
rect 1840 835 1890 850
rect 1940 1120 1990 1135
rect 1940 850 1955 1120
rect 1975 850 1990 1120
rect 1940 835 1990 850
rect 2040 1120 2090 1135
rect 2040 850 2055 1120
rect 2075 850 2090 1120
rect 2040 835 2090 850
rect 1410 820 1460 835
<< ndiffc >>
rect -325 425 -305 695
rect -225 425 -205 695
rect -125 425 -105 695
rect -25 425 -5 695
rect 75 425 95 695
rect 175 425 195 695
rect 305 425 325 695
rect 405 425 425 695
rect 485 425 505 695
rect 585 425 605 695
rect 685 425 705 695
rect 765 425 785 695
rect 865 425 885 695
rect 965 425 985 695
rect 1045 425 1065 695
rect 1145 425 1165 695
rect 1245 425 1265 695
rect 1325 425 1345 695
rect 1425 425 1445 695
rect 1555 410 1575 680
rect 1655 410 1675 680
rect 1755 410 1775 680
rect 1855 410 1875 680
rect 1955 410 1975 680
rect 2055 410 2075 680
rect -35 -25 -15 245
rect 65 -25 85 245
rect 165 -25 185 245
rect 265 -25 285 245
rect 365 -25 385 245
rect 465 -25 485 245
rect 565 -25 585 245
rect 665 -25 685 245
rect 765 -25 785 245
rect 865 -25 885 245
rect 965 -25 985 245
rect 1065 -25 1085 245
rect 1165 -25 1185 245
rect 1265 -25 1285 245
rect 1365 -25 1385 245
rect 1465 -25 1485 245
rect 1565 -25 1585 245
rect 1665 -25 1685 245
rect 1765 -25 1785 245
<< pdiffc >>
rect -35 1285 -15 1555
rect 65 1285 85 1555
rect 165 1285 185 1555
rect 265 1285 285 1555
rect 365 1285 385 1555
rect 465 1285 485 1555
rect 565 1285 585 1555
rect 665 1285 685 1555
rect 765 1285 785 1555
rect 865 1285 885 1555
rect 965 1285 985 1555
rect 1065 1285 1085 1555
rect 1165 1285 1185 1555
rect 1265 1285 1285 1555
rect 1365 1285 1385 1555
rect 1465 1285 1485 1555
rect 1565 1285 1585 1555
rect 1665 1285 1685 1555
rect 1765 1285 1785 1555
rect -725 835 -705 1105
rect -625 835 -605 1105
rect -525 835 -505 1105
rect -425 835 -405 1105
rect -325 835 -305 1105
rect -225 835 -205 1105
rect -125 835 -105 1105
rect -25 835 -5 1105
rect 75 835 95 1105
rect 175 835 195 1105
rect 305 835 325 1105
rect 405 835 425 1105
rect 485 835 505 1105
rect 585 835 605 1105
rect 685 835 705 1105
rect 765 835 785 1105
rect 865 835 885 1105
rect 965 835 985 1105
rect 1045 835 1065 1105
rect 1145 835 1165 1105
rect 1245 835 1265 1105
rect 1325 835 1345 1105
rect 1425 835 1445 1105
rect 1555 850 1575 1120
rect 1655 850 1675 1120
rect 1755 850 1775 1120
rect 1855 850 1875 1120
rect 1955 850 1975 1120
rect 2055 850 2075 1120
<< psubdiff >>
rect 240 695 290 710
rect 240 425 255 695
rect 275 425 290 695
rect 240 410 290 425
rect 1460 695 1510 710
rect 1460 425 1475 695
rect 1495 425 1510 695
rect 1460 410 1510 425
rect -340 245 -50 260
rect -340 -25 -325 245
rect -65 -25 -50 245
rect -340 -40 -50 -25
rect 1800 245 2090 260
rect 1800 -25 1815 245
rect 2075 -25 2090 245
rect 1800 -40 2090 -25
<< nsubdiff >>
rect -340 1555 -50 1570
rect -340 1285 -325 1555
rect -65 1285 -50 1555
rect -340 1270 -50 1285
rect 1800 1555 2090 1570
rect 1800 1285 1815 1555
rect 2075 1285 2090 1555
rect 1800 1270 2090 1285
rect 240 1105 290 1120
rect 240 835 255 1105
rect 275 835 290 1105
rect 240 820 290 835
rect 1460 1105 1510 1120
rect 1460 835 1475 1105
rect 1495 835 1510 1105
rect 1460 820 1510 835
<< psubdiffcont >>
rect 255 425 275 695
rect 1475 425 1495 695
rect -325 -25 -65 245
rect 1815 -25 2075 245
<< nsubdiffcont >>
rect -325 1285 -65 1555
rect 1815 1285 2075 1555
rect 255 835 275 1105
rect 1475 835 1495 1105
<< poly >>
rect 0 1570 50 1585
rect 100 1570 150 1585
rect 200 1570 250 1585
rect 300 1570 350 1585
rect 400 1570 450 1585
rect 500 1570 550 1585
rect 600 1570 650 1585
rect 700 1570 750 1585
rect 800 1570 850 1585
rect 900 1570 950 1585
rect 1000 1570 1050 1585
rect 1100 1570 1150 1585
rect 1200 1570 1250 1585
rect 1300 1570 1350 1585
rect 1400 1570 1450 1585
rect 1500 1570 1550 1585
rect 1600 1570 1650 1585
rect 1700 1570 1750 1585
rect 0 1245 50 1270
rect 0 1225 15 1245
rect 35 1225 50 1245
rect 0 1215 50 1225
rect 100 1245 150 1270
rect 100 1225 115 1245
rect 135 1225 150 1245
rect 100 1215 150 1225
rect 200 1245 250 1270
rect 200 1225 215 1245
rect 235 1225 250 1245
rect 200 1215 250 1225
rect 300 1245 350 1270
rect 300 1225 315 1245
rect 335 1225 350 1245
rect 300 1215 350 1225
rect 400 1245 450 1270
rect 400 1225 415 1245
rect 435 1225 450 1245
rect 400 1215 450 1225
rect 500 1245 550 1270
rect 500 1225 515 1245
rect 535 1225 550 1245
rect 500 1215 550 1225
rect 600 1245 650 1270
rect 600 1225 615 1245
rect 635 1225 650 1245
rect 600 1215 650 1225
rect 700 1245 750 1270
rect 700 1225 715 1245
rect 735 1225 750 1245
rect 700 1215 750 1225
rect 800 1245 850 1270
rect 800 1225 815 1245
rect 835 1225 850 1245
rect 800 1215 850 1225
rect 900 1245 950 1270
rect 900 1225 915 1245
rect 935 1225 950 1245
rect 900 1215 950 1225
rect 1000 1245 1050 1270
rect 1000 1225 1015 1245
rect 1035 1225 1050 1245
rect 1000 1215 1050 1225
rect 1100 1245 1150 1270
rect 1100 1225 1115 1245
rect 1135 1225 1150 1245
rect 1100 1215 1150 1225
rect 1200 1245 1250 1270
rect 1200 1225 1215 1245
rect 1235 1225 1250 1245
rect 1200 1215 1250 1225
rect 1300 1245 1350 1270
rect 1300 1225 1315 1245
rect 1335 1225 1350 1245
rect 1300 1215 1350 1225
rect 1400 1245 1450 1270
rect 1400 1225 1415 1245
rect 1435 1225 1450 1245
rect 1400 1215 1450 1225
rect 1500 1245 1550 1270
rect 1500 1225 1515 1245
rect 1535 1225 1550 1245
rect 1500 1215 1550 1225
rect 1600 1245 1650 1270
rect 1600 1225 1615 1245
rect 1635 1225 1650 1245
rect 1600 1215 1650 1225
rect 1700 1245 1750 1270
rect 1700 1225 1715 1245
rect 1735 1225 1750 1245
rect 1700 1215 1750 1225
rect 1990 1180 2040 1190
rect -690 1165 -640 1175
rect -690 1145 -675 1165
rect -655 1145 -640 1165
rect -690 1120 -640 1145
rect -590 1165 -540 1175
rect -590 1145 -575 1165
rect -555 1145 -540 1165
rect -590 1120 -540 1145
rect -490 1165 -440 1175
rect -490 1145 -475 1165
rect -455 1145 -440 1165
rect -490 1120 -440 1145
rect -390 1165 -340 1175
rect -390 1145 -375 1165
rect -355 1145 -340 1165
rect -390 1120 -340 1145
rect -290 1165 -240 1175
rect -290 1145 -275 1165
rect -255 1145 -240 1165
rect -290 1120 -240 1145
rect -190 1165 -140 1175
rect -190 1145 -175 1165
rect -155 1145 -140 1165
rect -190 1120 -140 1145
rect -90 1165 -40 1175
rect -90 1145 -75 1165
rect -55 1145 -40 1165
rect -90 1120 -40 1145
rect 10 1165 60 1175
rect 10 1145 25 1165
rect 45 1145 60 1165
rect 10 1120 60 1145
rect 110 1165 160 1175
rect 110 1145 125 1165
rect 145 1145 160 1165
rect 110 1120 160 1145
rect 210 1165 1410 1175
rect 210 1145 225 1165
rect 245 1145 1410 1165
rect 1990 1160 2005 1180
rect 2025 1160 2040 1180
rect 210 1135 1410 1145
rect 1590 1135 1640 1150
rect 1690 1135 1740 1150
rect 1790 1135 1840 1150
rect 1890 1135 1940 1150
rect 1990 1135 2040 1160
rect 340 1120 390 1135
rect 520 1120 570 1135
rect 620 1120 670 1135
rect 800 1120 850 1135
rect 900 1120 950 1135
rect 1080 1120 1130 1135
rect 1180 1120 1230 1135
rect 1360 1120 1410 1135
rect -690 805 -640 820
rect -590 805 -540 820
rect -490 805 -440 820
rect -390 805 -340 820
rect -290 805 -240 820
rect -190 805 -140 820
rect -90 805 -40 820
rect 10 805 60 820
rect 110 805 160 820
rect 340 805 390 820
rect 520 805 570 820
rect 620 805 670 820
rect 800 805 850 820
rect 900 805 950 820
rect 1080 805 1130 820
rect 1180 805 1230 820
rect 1360 805 1410 820
rect 1590 810 1640 835
rect 435 795 475 805
rect 1590 800 1605 810
rect 435 775 445 795
rect 465 775 475 795
rect 1510 790 1605 800
rect 1625 790 1640 810
rect 1510 780 1640 790
rect 1690 810 1740 835
rect 1690 790 1705 810
rect 1725 790 1740 810
rect 1690 780 1740 790
rect 1790 810 1840 835
rect 1790 790 1805 810
rect 1825 790 1840 810
rect 1790 780 1840 790
rect 1890 810 1940 835
rect 1990 820 2040 835
rect 1890 790 1905 810
rect 1925 790 1940 810
rect 1890 780 1940 790
rect 435 755 735 775
rect 1510 765 1530 780
rect 695 735 705 755
rect 725 735 735 755
rect 695 725 735 735
rect 1490 755 1530 765
rect 1490 735 1500 755
rect 1520 735 1530 755
rect 1490 725 1530 735
rect 1590 740 1640 750
rect -290 710 -240 725
rect -190 710 -140 725
rect -90 710 -40 725
rect 10 710 60 725
rect 110 710 160 725
rect 340 710 390 725
rect 520 710 570 725
rect 620 710 670 725
rect 800 710 850 725
rect 900 710 950 725
rect 1080 710 1130 725
rect 1180 710 1230 725
rect 1360 710 1410 725
rect 1590 720 1605 740
rect 1625 720 1640 740
rect 1590 695 1640 720
rect 1690 740 1740 750
rect 1690 720 1705 740
rect 1725 720 1740 740
rect 1690 695 1740 720
rect 1790 740 1840 750
rect 1790 720 1805 740
rect 1825 720 1840 740
rect 1790 695 1840 720
rect 1890 740 1940 750
rect 1890 720 1905 740
rect 1925 720 1940 740
rect 1890 695 1940 720
rect 1990 695 2040 710
rect -290 385 -240 410
rect -290 365 -275 385
rect -255 365 -240 385
rect -290 355 -240 365
rect -190 385 -140 410
rect -190 365 -175 385
rect -155 365 -140 385
rect -190 355 -140 365
rect -90 385 -40 410
rect -90 365 -75 385
rect -55 365 -40 385
rect -90 355 -40 365
rect 10 385 60 410
rect 10 365 25 385
rect 45 365 60 385
rect 10 355 60 365
rect 110 385 160 410
rect 340 395 390 410
rect 520 395 570 410
rect 620 395 670 410
rect 800 395 850 410
rect 900 395 950 410
rect 1080 395 1130 410
rect 1180 395 1230 410
rect 1360 395 1410 410
rect 110 365 125 385
rect 145 365 160 385
rect 110 355 160 365
rect 205 385 1410 395
rect 205 365 215 385
rect 235 365 1410 385
rect 1590 380 1640 395
rect 1690 380 1740 395
rect 1790 380 1840 395
rect 1890 380 1940 395
rect 205 355 1410 365
rect 1990 370 2040 395
rect 1990 350 2005 370
rect 2025 350 2040 370
rect 1990 340 2040 350
rect 0 305 50 315
rect 0 285 15 305
rect 35 285 50 305
rect 0 260 50 285
rect 100 305 150 315
rect 100 285 115 305
rect 135 285 150 305
rect 100 260 150 285
rect 200 305 250 315
rect 200 285 215 305
rect 235 285 250 305
rect 200 260 250 285
rect 300 305 350 315
rect 300 285 315 305
rect 335 285 350 305
rect 300 260 350 285
rect 400 305 450 315
rect 400 285 415 305
rect 435 285 450 305
rect 400 260 450 285
rect 500 305 550 315
rect 500 285 515 305
rect 535 285 550 305
rect 500 260 550 285
rect 600 305 650 315
rect 600 285 615 305
rect 635 285 650 305
rect 600 260 650 285
rect 700 305 750 315
rect 700 285 715 305
rect 735 285 750 305
rect 700 260 750 285
rect 800 305 850 315
rect 800 285 815 305
rect 835 285 850 305
rect 800 260 850 285
rect 900 305 950 315
rect 900 285 915 305
rect 935 285 950 305
rect 900 260 950 285
rect 1000 305 1050 315
rect 1000 285 1015 305
rect 1035 285 1050 305
rect 1000 260 1050 285
rect 1100 305 1150 315
rect 1100 285 1115 305
rect 1135 285 1150 305
rect 1100 260 1150 285
rect 1200 305 1250 315
rect 1200 285 1215 305
rect 1235 285 1250 305
rect 1200 260 1250 285
rect 1300 305 1350 315
rect 1300 285 1315 305
rect 1335 285 1350 305
rect 1300 260 1350 285
rect 1400 305 1450 315
rect 1400 285 1415 305
rect 1435 285 1450 305
rect 1400 260 1450 285
rect 1500 305 1550 315
rect 1500 285 1515 305
rect 1535 285 1550 305
rect 1500 260 1550 285
rect 1600 305 1650 315
rect 1600 285 1615 305
rect 1635 285 1650 305
rect 1600 260 1650 285
rect 1700 305 1750 315
rect 1700 285 1715 305
rect 1735 285 1750 305
rect 1700 260 1750 285
rect 0 -55 50 -40
rect 100 -55 150 -40
rect 200 -55 250 -40
rect 300 -55 350 -40
rect 400 -55 450 -40
rect 500 -55 550 -40
rect 600 -55 650 -40
rect 700 -55 750 -40
rect 800 -55 850 -40
rect 900 -55 950 -40
rect 1000 -55 1050 -40
rect 1100 -55 1150 -40
rect 1200 -55 1250 -40
rect 1300 -55 1350 -40
rect 1400 -55 1450 -40
rect 1500 -55 1550 -40
rect 1600 -55 1650 -40
rect 1700 -55 1750 -40
<< polycont >>
rect 15 1225 35 1245
rect 115 1225 135 1245
rect 215 1225 235 1245
rect 315 1225 335 1245
rect 415 1225 435 1245
rect 515 1225 535 1245
rect 615 1225 635 1245
rect 715 1225 735 1245
rect 815 1225 835 1245
rect 915 1225 935 1245
rect 1015 1225 1035 1245
rect 1115 1225 1135 1245
rect 1215 1225 1235 1245
rect 1315 1225 1335 1245
rect 1415 1225 1435 1245
rect 1515 1225 1535 1245
rect 1615 1225 1635 1245
rect 1715 1225 1735 1245
rect -675 1145 -655 1165
rect -575 1145 -555 1165
rect -475 1145 -455 1165
rect -375 1145 -355 1165
rect -275 1145 -255 1165
rect -175 1145 -155 1165
rect -75 1145 -55 1165
rect 25 1145 45 1165
rect 125 1145 145 1165
rect 225 1145 245 1165
rect 2005 1160 2025 1180
rect 445 775 465 795
rect 1605 790 1625 810
rect 1705 790 1725 810
rect 1805 790 1825 810
rect 1905 790 1925 810
rect 705 735 725 755
rect 1500 735 1520 755
rect 1605 720 1625 740
rect 1705 720 1725 740
rect 1805 720 1825 740
rect 1905 720 1925 740
rect -275 365 -255 385
rect -175 365 -155 385
rect -75 365 -55 385
rect 25 365 45 385
rect 125 365 145 385
rect 215 365 235 385
rect 2005 350 2025 370
rect 15 285 35 305
rect 115 285 135 305
rect 215 285 235 305
rect 315 285 335 305
rect 415 285 435 305
rect 515 285 535 305
rect 615 285 635 305
rect 715 285 735 305
rect 815 285 835 305
rect 915 285 935 305
rect 1015 285 1035 305
rect 1115 285 1135 305
rect 1215 285 1235 305
rect 1315 285 1335 305
rect 1415 285 1435 305
rect 1515 285 1535 305
rect 1615 285 1635 305
rect 1715 285 1735 305
<< locali >>
rect 65 1585 1685 1605
rect 65 1565 85 1585
rect 265 1565 285 1585
rect 465 1565 485 1585
rect 665 1565 685 1585
rect 865 1565 885 1585
rect 1065 1565 1085 1585
rect 1265 1565 1285 1585
rect 1465 1565 1485 1585
rect 1665 1565 1685 1585
rect -335 1555 -5 1565
rect -335 1285 -325 1555
rect -65 1285 -35 1555
rect -15 1285 -5 1555
rect -335 1275 -5 1285
rect 55 1555 95 1565
rect 55 1285 65 1555
rect 85 1285 95 1555
rect 55 1275 95 1285
rect 155 1555 195 1565
rect 155 1285 165 1555
rect 185 1285 195 1555
rect 155 1275 195 1285
rect 255 1555 295 1565
rect 255 1285 265 1555
rect 285 1285 295 1555
rect 255 1275 295 1285
rect 355 1555 395 1565
rect 355 1285 365 1555
rect 385 1285 395 1555
rect 355 1275 395 1285
rect 455 1555 495 1565
rect 455 1285 465 1555
rect 485 1285 495 1555
rect 455 1275 495 1285
rect 555 1555 595 1565
rect 555 1285 565 1555
rect 585 1285 595 1555
rect 555 1275 595 1285
rect 655 1555 695 1565
rect 655 1285 665 1555
rect 685 1285 695 1555
rect 655 1275 695 1285
rect 755 1555 795 1565
rect 755 1285 765 1555
rect 785 1285 795 1555
rect 755 1275 795 1285
rect 855 1555 895 1565
rect 855 1285 865 1555
rect 885 1285 895 1555
rect 855 1275 895 1285
rect 955 1555 995 1565
rect 955 1285 965 1555
rect 985 1285 995 1555
rect 955 1275 995 1285
rect 1055 1555 1095 1565
rect 1055 1285 1065 1555
rect 1085 1285 1095 1555
rect 1055 1275 1095 1285
rect 1155 1555 1195 1565
rect 1155 1285 1165 1555
rect 1185 1285 1195 1555
rect 1155 1275 1195 1285
rect 1255 1555 1295 1565
rect 1255 1285 1265 1555
rect 1285 1285 1295 1555
rect 1255 1275 1295 1285
rect 1355 1555 1395 1565
rect 1355 1285 1365 1555
rect 1385 1285 1395 1555
rect 1355 1275 1395 1285
rect 1455 1555 1495 1565
rect 1455 1285 1465 1555
rect 1485 1285 1495 1555
rect 1455 1275 1495 1285
rect 1555 1555 1595 1565
rect 1555 1285 1565 1555
rect 1585 1285 1595 1555
rect 1555 1275 1595 1285
rect 1655 1555 1695 1565
rect 1655 1285 1665 1555
rect 1685 1285 1695 1555
rect 1655 1275 1695 1285
rect 1755 1555 2085 1565
rect 1755 1285 1765 1555
rect 1785 1285 1815 1555
rect 2075 1285 2085 1555
rect 1755 1275 2085 1285
rect -45 1255 -5 1275
rect 165 1255 185 1275
rect 365 1255 385 1275
rect 765 1255 785 1275
rect 965 1255 985 1275
rect 1365 1255 1385 1275
rect 1565 1255 1585 1275
rect 1755 1255 1795 1275
rect -45 1245 50 1255
rect -45 1225 15 1245
rect 35 1225 50 1245
rect -45 1215 50 1225
rect 100 1245 1650 1255
rect 100 1225 115 1245
rect 135 1225 215 1245
rect 235 1225 315 1245
rect 335 1225 415 1245
rect 435 1225 515 1245
rect 535 1225 615 1245
rect 635 1225 715 1245
rect 735 1225 815 1245
rect 835 1225 915 1245
rect 935 1225 1015 1245
rect 1035 1225 1115 1245
rect 1135 1225 1215 1245
rect 1235 1225 1315 1245
rect 1335 1225 1415 1245
rect 1435 1225 1515 1245
rect 1535 1225 1615 1245
rect 1635 1225 1650 1245
rect 100 1215 1650 1225
rect 1700 1245 1795 1255
rect 1700 1225 1715 1245
rect 1735 1225 1795 1245
rect 1700 1215 1795 1225
rect -735 1165 -640 1175
rect -735 1145 -675 1165
rect -655 1145 -640 1165
rect -735 1135 -640 1145
rect -615 1165 260 1175
rect -615 1145 -575 1165
rect -555 1145 -475 1165
rect -455 1145 -375 1165
rect -355 1145 -275 1165
rect -255 1145 -175 1165
rect -155 1145 -75 1165
rect -55 1145 25 1165
rect 45 1145 125 1165
rect 145 1145 225 1165
rect 245 1145 260 1165
rect -615 1135 260 1145
rect -735 1105 -695 1135
rect -615 1115 -595 1135
rect -225 1115 -205 1135
rect 175 1115 195 1135
rect -735 835 -725 1105
rect -705 835 -695 1105
rect -735 825 -695 835
rect -635 1105 -595 1115
rect -635 835 -625 1105
rect -605 835 -595 1105
rect -635 825 -595 835
rect -535 1105 -495 1115
rect -535 835 -525 1105
rect -505 835 -495 1105
rect -535 825 -495 835
rect -435 1105 -395 1115
rect -435 835 -425 1105
rect -405 835 -395 1105
rect -435 825 -395 835
rect -335 1105 -295 1115
rect -335 835 -325 1105
rect -305 835 -295 1105
rect -335 825 -295 835
rect -235 1105 -195 1115
rect -235 835 -225 1105
rect -205 835 -195 1105
rect -235 825 -195 835
rect -135 1105 -95 1115
rect -135 835 -125 1105
rect -105 835 -95 1105
rect -135 825 -95 835
rect -35 1105 5 1115
rect -35 835 -25 1105
rect -5 835 5 1105
rect -35 825 5 835
rect 65 1105 105 1115
rect 65 835 75 1105
rect 95 835 105 1105
rect 65 825 105 835
rect 165 1105 205 1115
rect 165 835 175 1105
rect 195 835 205 1105
rect -635 805 -615 825
rect -740 785 -615 805
rect -425 805 -405 825
rect -25 805 -5 825
rect -425 785 -5 805
rect -25 780 -5 785
rect 165 800 205 835
rect 245 1105 335 1115
rect 245 835 255 1105
rect 275 835 305 1105
rect 325 835 335 1105
rect 245 825 335 835
rect 165 780 175 800
rect 195 780 205 800
rect 355 805 375 1215
rect 415 1175 1435 1195
rect 415 1115 435 1175
rect 495 1135 1055 1155
rect 495 1115 515 1135
rect 1035 1115 1055 1135
rect 1415 1115 1435 1175
rect 1990 1180 2085 1190
rect 1555 1150 1965 1170
rect 1990 1160 2005 1180
rect 2025 1160 2085 1180
rect 1990 1150 2085 1160
rect 1555 1130 1575 1150
rect 1755 1130 1775 1150
rect 1945 1130 1965 1150
rect 1545 1120 1585 1130
rect 395 1105 435 1115
rect 395 835 405 1105
rect 425 835 435 1105
rect 395 825 435 835
rect 475 1105 515 1115
rect 475 835 485 1105
rect 505 835 515 1105
rect 475 825 515 835
rect 575 1105 615 1115
rect 575 835 585 1105
rect 605 835 615 1105
rect 575 825 615 835
rect 675 1105 715 1115
rect 675 835 685 1105
rect 705 835 715 1105
rect 675 825 715 835
rect 755 1105 795 1115
rect 755 835 765 1105
rect 785 835 795 1105
rect 755 825 795 835
rect 855 1105 895 1115
rect 855 835 865 1105
rect 885 835 895 1105
rect 855 825 895 835
rect 955 1105 995 1115
rect 955 835 965 1105
rect 985 835 995 1105
rect 955 825 995 835
rect 1035 1105 1075 1115
rect 1035 835 1045 1105
rect 1065 835 1075 1105
rect 1035 825 1075 835
rect 1135 1105 1175 1115
rect 1135 835 1145 1105
rect 1165 835 1175 1105
rect 1135 825 1175 835
rect 1235 1105 1275 1115
rect 1235 835 1245 1105
rect 1265 835 1275 1105
rect 1235 825 1275 835
rect 1315 1105 1355 1115
rect 1315 835 1325 1105
rect 1345 835 1355 1105
rect 1315 825 1355 835
rect 1415 1105 1505 1115
rect 1415 835 1425 1105
rect 1445 835 1475 1105
rect 1495 835 1505 1105
rect 1545 850 1555 1120
rect 1575 850 1585 1120
rect 1545 840 1585 850
rect 1645 1120 1685 1130
rect 1645 850 1655 1120
rect 1675 850 1685 1120
rect 1645 840 1685 850
rect 1745 1120 1785 1130
rect 1745 850 1755 1120
rect 1775 850 1785 1120
rect 1745 840 1785 850
rect 1845 1120 1885 1130
rect 1845 850 1855 1120
rect 1875 850 1885 1120
rect 1845 840 1885 850
rect 1945 1120 1985 1130
rect 1945 850 1955 1120
rect 1975 850 1985 1120
rect 1945 840 1985 850
rect 2045 1120 2085 1150
rect 2045 850 2055 1120
rect 2075 850 2085 1120
rect 2045 840 2085 850
rect 1415 825 1505 835
rect 655 805 695 825
rect 765 805 785 825
rect 965 805 985 825
rect 1315 805 1335 825
rect 1655 820 1675 840
rect 1855 820 1875 840
rect 1590 810 2090 820
rect 355 795 475 805
rect 355 785 445 795
rect -25 770 15 780
rect 165 770 205 780
rect 435 775 445 785
rect 465 775 475 795
rect -25 750 -15 770
rect 5 750 15 770
rect 435 765 475 775
rect -25 740 15 750
rect 655 745 675 805
rect 765 785 1570 805
rect -25 705 -5 740
rect 355 725 675 745
rect 695 755 735 765
rect 695 735 705 755
rect 725 735 735 755
rect 1490 755 1530 765
rect 1490 745 1500 755
rect 695 725 735 735
rect 765 735 1500 745
rect 1520 735 1530 755
rect 765 725 1530 735
rect 1550 750 1570 785
rect 1590 790 1605 810
rect 1625 790 1705 810
rect 1725 790 1805 810
rect 1825 790 1905 810
rect 1925 800 2090 810
rect 1925 790 1940 800
rect 1590 780 1940 790
rect 1550 740 1940 750
rect 1550 730 1605 740
rect -335 695 -295 705
rect -335 425 -325 695
rect -305 425 -295 695
rect -335 395 -295 425
rect -235 695 -195 705
rect -235 425 -225 695
rect -205 425 -195 695
rect -235 415 -195 425
rect -135 695 -95 705
rect -135 425 -125 695
rect -105 425 -95 695
rect -135 415 -95 425
rect -35 695 5 705
rect -35 425 -25 695
rect -5 425 5 695
rect -35 415 5 425
rect 65 695 105 705
rect 65 425 75 695
rect 95 425 105 695
rect 65 415 105 425
rect 165 695 205 705
rect 165 425 175 695
rect 195 425 205 695
rect 165 415 205 425
rect 245 695 335 705
rect 245 425 255 695
rect 275 425 305 695
rect 325 425 335 695
rect 245 415 335 425
rect -215 395 -195 415
rect -25 395 -5 415
rect 175 395 195 415
rect -335 385 -240 395
rect -335 365 -275 385
rect -255 365 -240 385
rect -335 355 -240 365
rect -215 385 245 395
rect -215 365 -175 385
rect -155 365 -75 385
rect -55 365 25 385
rect 45 365 125 385
rect 145 365 215 385
rect 235 365 245 385
rect -215 355 245 365
rect 355 315 375 725
rect 695 705 715 725
rect 765 705 785 725
rect 965 705 985 725
rect 1315 705 1335 725
rect 1590 720 1605 730
rect 1625 720 1705 740
rect 1725 720 1805 740
rect 1825 720 1905 740
rect 1925 730 1940 740
rect 1925 720 2090 730
rect 1590 710 2090 720
rect 395 695 435 705
rect 395 425 405 695
rect 425 425 435 695
rect 395 415 435 425
rect 475 695 515 705
rect 475 425 485 695
rect 505 425 515 695
rect 475 415 515 425
rect 575 695 615 705
rect 575 425 585 695
rect 605 425 615 695
rect 575 415 615 425
rect 675 695 715 705
rect 675 425 685 695
rect 705 425 715 695
rect 675 415 715 425
rect 755 695 795 705
rect 755 425 765 695
rect 785 425 795 695
rect 755 415 795 425
rect 855 695 895 705
rect 855 425 865 695
rect 885 425 895 695
rect 855 415 895 425
rect 955 695 995 705
rect 955 425 965 695
rect 985 425 995 695
rect 955 415 995 425
rect 1035 695 1075 705
rect 1035 425 1045 695
rect 1065 425 1075 695
rect 1035 415 1075 425
rect 1135 695 1175 705
rect 1135 425 1145 695
rect 1165 425 1175 695
rect 1135 415 1175 425
rect 1235 695 1275 705
rect 1235 425 1245 695
rect 1265 425 1275 695
rect 1235 415 1275 425
rect 1315 695 1355 705
rect 1315 425 1325 695
rect 1345 425 1355 695
rect 1315 415 1355 425
rect 1415 695 1505 705
rect 1415 425 1425 695
rect 1445 425 1475 695
rect 1495 425 1505 695
rect 1655 690 1675 710
rect 1855 690 1875 710
rect 1415 415 1505 425
rect 1545 680 1585 690
rect 415 355 435 415
rect 495 395 515 415
rect 1035 395 1055 415
rect 495 375 1055 395
rect 1415 355 1435 415
rect 1545 410 1555 680
rect 1575 410 1585 680
rect 1545 400 1585 410
rect 1645 680 1685 690
rect 1645 410 1655 680
rect 1675 410 1685 680
rect 1645 400 1685 410
rect 1745 680 1785 690
rect 1745 410 1755 680
rect 1775 410 1785 680
rect 1745 400 1785 410
rect 1845 680 1885 690
rect 1845 410 1855 680
rect 1875 410 1885 680
rect 1845 400 1885 410
rect 1945 680 1985 690
rect 1945 410 1955 680
rect 1975 410 1985 680
rect 1945 400 1985 410
rect 2045 680 2085 690
rect 2045 410 2055 680
rect 2075 410 2085 680
rect 1555 380 1575 400
rect 1755 380 1775 400
rect 1945 380 1965 400
rect 2045 380 2085 410
rect 1555 360 1965 380
rect 1990 370 2085 380
rect 415 335 1435 355
rect 1990 350 2005 370
rect 2025 350 2085 370
rect 1990 340 2085 350
rect -45 305 50 315
rect -45 285 15 305
rect 35 285 50 305
rect -45 275 50 285
rect 100 305 1650 315
rect 100 285 115 305
rect 135 285 215 305
rect 235 285 315 305
rect 335 285 415 305
rect 435 285 515 305
rect 535 285 615 305
rect 635 285 715 305
rect 735 285 815 305
rect 835 285 915 305
rect 935 285 1015 305
rect 1035 285 1115 305
rect 1135 285 1215 305
rect 1235 285 1315 305
rect 1335 285 1415 305
rect 1435 285 1515 305
rect 1535 285 1615 305
rect 1635 285 1650 305
rect 100 275 1650 285
rect 1700 305 1795 315
rect 1700 285 1715 305
rect 1735 285 1795 305
rect 1700 275 1795 285
rect -45 255 -5 275
rect 165 255 185 275
rect 365 255 385 275
rect 765 255 785 275
rect 965 255 985 275
rect 1365 255 1385 275
rect 1565 255 1585 275
rect 1755 255 1795 275
rect -335 245 -5 255
rect -335 -25 -325 245
rect -65 -25 -35 245
rect -15 -25 -5 245
rect -335 -35 -5 -25
rect 55 245 95 255
rect 55 -25 65 245
rect 85 -25 95 245
rect 55 -35 95 -25
rect 155 245 195 255
rect 155 -25 165 245
rect 185 -25 195 245
rect 155 -35 195 -25
rect 255 245 295 255
rect 255 -25 265 245
rect 285 -25 295 245
rect 255 -35 295 -25
rect 355 245 395 255
rect 355 -25 365 245
rect 385 -25 395 245
rect 355 -35 395 -25
rect 455 245 495 255
rect 455 -25 465 245
rect 485 -25 495 245
rect 455 -35 495 -25
rect 555 245 595 255
rect 555 -25 565 245
rect 585 -25 595 245
rect 555 -35 595 -25
rect 655 245 695 255
rect 655 -25 665 245
rect 685 -25 695 245
rect 655 -35 695 -25
rect 755 245 795 255
rect 755 -25 765 245
rect 785 -25 795 245
rect 755 -35 795 -25
rect 855 245 895 255
rect 855 -25 865 245
rect 885 -25 895 245
rect 855 -35 895 -25
rect 955 245 995 255
rect 955 -25 965 245
rect 985 -25 995 245
rect 955 -35 995 -25
rect 1055 245 1095 255
rect 1055 -25 1065 245
rect 1085 -25 1095 245
rect 1055 -35 1095 -25
rect 1155 245 1195 255
rect 1155 -25 1165 245
rect 1185 -25 1195 245
rect 1155 -35 1195 -25
rect 1255 245 1295 255
rect 1255 -25 1265 245
rect 1285 -25 1295 245
rect 1255 -35 1295 -25
rect 1355 245 1395 255
rect 1355 -25 1365 245
rect 1385 -25 1395 245
rect 1355 -35 1395 -25
rect 1455 245 1495 255
rect 1455 -25 1465 245
rect 1485 -25 1495 245
rect 1455 -35 1495 -25
rect 1555 245 1595 255
rect 1555 -25 1565 245
rect 1585 -25 1595 245
rect 1555 -35 1595 -25
rect 1655 245 1695 255
rect 1655 -25 1665 245
rect 1685 -25 1695 245
rect 1655 -35 1695 -25
rect 1755 245 2085 255
rect 1755 -25 1765 245
rect 1785 -25 1815 245
rect 2075 -25 2085 245
rect 1755 -35 2085 -25
rect 65 -55 85 -35
rect 265 -55 285 -35
rect 465 -55 485 -35
rect 665 -55 685 -35
rect 865 -55 885 -35
rect 1065 -55 1085 -35
rect 1265 -55 1285 -35
rect 1465 -55 1485 -35
rect 1665 -55 1685 -35
rect 65 -75 1685 -55
<< viali >>
rect -325 1285 -65 1555
rect -35 1285 -15 1555
rect 565 1285 585 1555
rect 1165 1285 1185 1555
rect 1765 1285 1785 1555
rect 1815 1285 2075 1555
rect -725 835 -705 1105
rect -525 835 -505 1105
rect -325 835 -305 1105
rect -125 835 -105 1105
rect 75 835 95 1105
rect 255 835 275 1105
rect 305 835 325 1105
rect 175 780 195 800
rect 865 835 885 1105
rect 1245 835 1265 1105
rect 1425 835 1445 1105
rect 1475 835 1495 1105
rect 2055 850 2075 1120
rect -15 750 5 770
rect -325 425 -305 695
rect -125 425 -105 695
rect 75 425 95 695
rect 255 425 275 695
rect 305 425 325 695
rect 865 425 885 695
rect 1245 425 1265 695
rect 1425 425 1445 695
rect 1475 425 1495 695
rect 2055 410 2075 680
rect -325 -25 -65 245
rect -35 -25 -15 245
rect 565 -25 585 245
rect 1165 -25 1185 245
rect 1765 -25 1785 245
rect 1815 -25 2075 245
<< metal1 >>
rect -740 1555 2090 1570
rect -740 1285 -325 1555
rect -65 1285 -35 1555
rect -15 1285 565 1555
rect 585 1285 1165 1555
rect 1185 1285 1765 1555
rect 1785 1285 1815 1555
rect 2075 1285 2090 1555
rect -740 1120 2090 1285
rect -740 1105 2055 1120
rect -740 835 -725 1105
rect -705 835 -525 1105
rect -505 835 -325 1105
rect -305 835 -125 1105
rect -105 835 75 1105
rect 95 840 255 1105
rect 95 835 135 840
rect -740 820 135 835
rect 235 835 255 840
rect 275 835 305 1105
rect 325 835 865 1105
rect 885 835 1245 1105
rect 1265 835 1425 1105
rect 1445 835 1475 1105
rect 1495 850 2055 1105
rect 2075 850 2090 1120
rect 1495 835 2090 850
rect 235 820 2090 835
rect 165 800 205 810
rect 165 780 175 800
rect 195 785 205 800
rect 195 780 2090 785
rect -25 770 15 780
rect 165 770 2090 780
rect -25 750 -15 770
rect 5 755 15 770
rect 5 750 2090 755
rect -25 740 2090 750
rect -740 695 2090 710
rect -740 425 -325 695
rect -305 425 -125 695
rect -105 425 75 695
rect 95 425 255 695
rect 275 425 305 695
rect 325 425 865 695
rect 885 425 1245 695
rect 1265 425 1425 695
rect 1445 425 1475 695
rect 1495 680 2090 695
rect 1495 425 2055 680
rect -740 410 2055 425
rect 2075 410 2090 680
rect -740 245 2090 410
rect -740 -25 -325 245
rect -65 -25 -35 245
rect -15 -25 565 245
rect 585 -25 1165 245
rect 1185 -25 1765 245
rect 1785 -25 1815 245
rect 2075 -25 2090 245
rect -740 -40 2090 -25
<< labels >>
flabel metal1 2090 750 2090 750 3 FreeSans 160 0 0 0 Vb
port 1 e
flabel locali 2090 720 2090 720 3 FreeSans 160 0 0 0 Vcn
port 2 e
flabel locali 2090 810 2090 810 3 FreeSans 160 0 0 0 Vcp
port 3 e
flabel metal1 2090 775 2090 775 3 FreeSans 160 0 0 0 Vbp
port 4 e
flabel metal1 -740 1175 -740 1175 7 FreeSans 160 0 0 0 VP
port 5 w
flabel metal1 -740 355 -740 355 7 FreeSans 160 0 0 0 VN
port 6 w
<< end >>
