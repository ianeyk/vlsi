** SHIFT_REGISTER_INVERTER flat netlist
*--------BEGIN_X5->INVERTER
*.IOPIN VP
*.IOPIN VN
*.IPIN A
*.OPIN Y
*--------BEGIN_X5_XM1->SKY130_FD_PR__NFET_01V8
XM1_X5 DBAR1 A GND GND  SKY130_FD_PR__NFET_01V8 L=0.15 W=1 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___X5_XM1->SKY130_FD_PR__NFET_01V8
*--------BEGIN_X5_XM2->SKY130_FD_PR__PFET_01V8
XM2_X5 DBAR1 A VDD VDD  SKY130_FD_PR__PFET_01V8 L=0.15 W=4 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___X5_XM2->SKY130_FD_PR__PFET_01V8
*--------END___X5->INVERTER
*--------BEGIN_X6->INVERTER
*.IOPIN VP
*.IOPIN VN
*.IPIN A
*.OPIN Y
*--------BEGIN_X6_XM1->SKY130_FD_PR__NFET_01V8
XM1_X6 D1 DBAR1 GND GND  SKY130_FD_PR__NFET_01V8 L=0.15 W=1 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___X6_XM1->SKY130_FD_PR__NFET_01V8
*--------BEGIN_X6_XM2->SKY130_FD_PR__PFET_01V8
XM2_X6 D1 DBAR1 VDD VDD  SKY130_FD_PR__PFET_01V8 L=0.15 W=4 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___X6_XM2->SKY130_FD_PR__PFET_01V8
*--------END___X6->INVERTER
.end
