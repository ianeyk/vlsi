magic
tech sky130A
timestamp 1697031584
<< error_p >>
rect 125 2097 145 2100
rect 125 1833 128 2097
rect 142 1833 145 2097
rect 125 1830 145 1833
rect 325 2097 345 2100
rect 325 1833 328 2097
rect 342 1833 345 2097
rect 325 1830 345 1833
rect 525 2097 545 2100
rect 525 1833 528 2097
rect 542 1833 545 2097
rect 525 1830 545 1833
rect 725 2097 745 2100
rect 725 1833 728 2097
rect 742 1833 745 2097
rect 725 1830 745 1833
rect 925 2097 945 2100
rect 925 1833 928 2097
rect 942 1833 945 2097
rect 925 1830 945 1833
rect 1125 2097 1145 2100
rect 1125 1833 1128 2097
rect 1142 1833 1145 2097
rect 1125 1830 1145 1833
rect 125 1627 145 1630
rect 125 1363 128 1627
rect 142 1363 145 1627
rect 125 1360 145 1363
rect 1125 1627 1145 1630
rect 1125 1363 1128 1627
rect 1142 1363 1145 1627
rect 1125 1360 1145 1363
rect 125 1122 145 1125
rect 125 858 128 1122
rect 142 858 145 1122
rect 125 855 145 858
rect 325 1122 345 1125
rect 325 858 328 1122
rect 342 858 345 1122
rect 325 855 345 858
rect 525 1122 545 1125
rect 525 858 528 1122
rect 542 858 545 1122
rect 525 855 545 858
rect 725 1122 745 1125
rect 725 858 728 1122
rect 742 858 745 1122
rect 725 855 745 858
rect 925 1122 945 1125
rect 925 858 928 1122
rect 942 858 945 1122
rect 925 855 945 858
rect 1125 1122 1145 1125
rect 1125 858 1128 1122
rect 1142 858 1145 1122
rect 1125 855 1145 858
rect 125 -123 145 -120
rect 125 -387 128 -123
rect 142 -387 145 -123
rect 125 -390 145 -387
rect 325 -123 345 -120
rect 325 -387 328 -123
rect 342 -387 345 -123
rect 325 -390 345 -387
rect 525 -123 545 -120
rect 525 -387 528 -123
rect 542 -387 545 -123
rect 525 -390 545 -387
rect 725 -123 745 -120
rect 725 -387 728 -123
rect 742 -387 745 -123
rect 725 -390 745 -387
rect 925 -123 945 -120
rect 925 -387 928 -123
rect 942 -387 945 -123
rect 925 -390 945 -387
rect 1125 -123 1145 -120
rect 1125 -387 1128 -123
rect 1142 -387 1145 -123
rect 1125 -390 1145 -387
<< nwell >>
rect 90 775 1180 1160
rect -70 375 1340 775
<< nmos >>
rect 160 1815 210 2115
rect 260 1815 310 2115
rect 360 1815 410 2115
rect 460 1815 510 2115
rect 560 1815 610 2115
rect 660 1815 710 2115
rect 760 1815 810 2115
rect 860 1815 910 2115
rect 960 1815 1010 2115
rect 1060 1815 1110 2115
rect 160 1345 210 1645
rect 260 1345 310 1645
rect 360 1345 410 1645
rect 460 1345 510 1645
rect 560 1345 610 1645
rect 660 1345 710 1645
rect 760 1345 810 1645
rect 860 1345 910 1645
rect 960 1345 1010 1645
rect 1060 1345 1110 1645
rect 0 0 50 300
rect 100 0 150 300
rect 280 0 330 300
rect 380 0 430 300
rect 560 0 610 300
rect 660 0 710 300
rect 840 0 890 300
rect 940 0 990 300
rect 1120 0 1170 300
rect 1220 0 1270 300
rect 160 -405 210 -105
rect 260 -405 310 -105
rect 360 -405 410 -105
rect 460 -405 510 -105
rect 560 -405 610 -105
rect 660 -405 710 -105
rect 760 -405 810 -105
rect 860 -405 910 -105
rect 960 -405 1010 -105
rect 1060 -405 1110 -105
<< pmos >>
rect 160 840 210 1140
rect 260 840 310 1140
rect 360 840 410 1140
rect 460 840 510 1140
rect 560 840 610 1140
rect 660 840 710 1140
rect 760 840 810 1140
rect 860 840 910 1140
rect 960 840 1010 1140
rect 1060 840 1110 1140
rect 0 395 50 695
rect 100 395 150 695
rect 280 395 330 695
rect 380 395 430 695
rect 560 395 610 695
rect 660 395 710 695
rect 840 395 890 695
rect 940 395 990 695
rect 1120 395 1170 695
rect 1220 395 1270 695
<< ndiff >>
rect 110 2100 160 2115
rect 110 1830 125 2100
rect 145 1830 160 2100
rect 110 1815 160 1830
rect 210 2100 260 2115
rect 210 1830 225 2100
rect 245 1830 260 2100
rect 210 1815 260 1830
rect 310 2100 360 2115
rect 310 1830 325 2100
rect 345 1830 360 2100
rect 310 1815 360 1830
rect 410 2100 460 2115
rect 410 1830 425 2100
rect 445 1830 460 2100
rect 410 1815 460 1830
rect 510 2100 560 2115
rect 510 1830 525 2100
rect 545 1830 560 2100
rect 510 1815 560 1830
rect 610 2100 660 2115
rect 610 1830 625 2100
rect 645 1830 660 2100
rect 610 1815 660 1830
rect 710 2100 760 2115
rect 710 1830 725 2100
rect 745 1830 760 2100
rect 710 1815 760 1830
rect 810 2100 860 2115
rect 810 1830 825 2100
rect 845 1830 860 2100
rect 810 1815 860 1830
rect 910 2100 960 2115
rect 910 1830 925 2100
rect 945 1830 960 2100
rect 910 1815 960 1830
rect 1010 2100 1060 2115
rect 1010 1830 1025 2100
rect 1045 1830 1060 2100
rect 1010 1815 1060 1830
rect 1110 2100 1160 2115
rect 1110 1830 1125 2100
rect 1145 1830 1160 2100
rect 1110 1815 1160 1830
rect 110 1630 160 1645
rect 110 1360 125 1630
rect 145 1360 160 1630
rect 110 1345 160 1360
rect 210 1630 260 1645
rect 210 1360 225 1630
rect 245 1360 260 1630
rect 210 1345 260 1360
rect 310 1630 360 1645
rect 310 1360 325 1630
rect 345 1360 360 1630
rect 310 1345 360 1360
rect 410 1630 460 1645
rect 410 1360 425 1630
rect 445 1360 460 1630
rect 410 1345 460 1360
rect 510 1630 560 1645
rect 510 1360 525 1630
rect 545 1360 560 1630
rect 510 1345 560 1360
rect 610 1630 660 1645
rect 610 1360 625 1630
rect 645 1360 660 1630
rect 610 1345 660 1360
rect 710 1630 760 1645
rect 710 1360 725 1630
rect 745 1360 760 1630
rect 710 1345 760 1360
rect 810 1630 860 1645
rect 810 1360 825 1630
rect 845 1360 860 1630
rect 810 1345 860 1360
rect 910 1630 960 1645
rect 910 1360 925 1630
rect 945 1360 960 1630
rect 910 1345 960 1360
rect 1010 1630 1060 1645
rect 1010 1360 1025 1630
rect 1045 1360 1060 1630
rect 1010 1345 1060 1360
rect 1110 1630 1160 1645
rect 1110 1360 1125 1630
rect 1145 1360 1160 1630
rect 1110 1345 1160 1360
rect -50 285 0 300
rect -50 15 -35 285
rect -15 15 0 285
rect -50 0 0 15
rect 50 285 100 300
rect 50 15 65 285
rect 85 15 100 285
rect 50 0 100 15
rect 150 285 200 300
rect 150 15 165 285
rect 185 15 200 285
rect 150 0 200 15
rect 230 285 280 300
rect 230 15 245 285
rect 265 15 280 285
rect 230 0 280 15
rect 330 285 380 300
rect 330 15 345 285
rect 365 15 380 285
rect 330 0 380 15
rect 430 285 480 300
rect 430 15 445 285
rect 465 15 480 285
rect 430 0 480 15
rect 510 285 560 300
rect 510 15 525 285
rect 545 15 560 285
rect 510 0 560 15
rect 610 285 660 300
rect 610 15 625 285
rect 645 15 660 285
rect 610 0 660 15
rect 710 285 760 300
rect 710 15 725 285
rect 745 15 760 285
rect 710 0 760 15
rect 790 285 840 300
rect 790 15 805 285
rect 825 15 840 285
rect 790 0 840 15
rect 890 285 940 300
rect 890 15 905 285
rect 925 15 940 285
rect 890 0 940 15
rect 990 285 1040 300
rect 990 15 1005 285
rect 1025 15 1040 285
rect 990 0 1040 15
rect 1070 285 1120 300
rect 1070 15 1085 285
rect 1105 15 1120 285
rect 1070 0 1120 15
rect 1170 285 1220 300
rect 1170 15 1185 285
rect 1205 15 1220 285
rect 1170 0 1220 15
rect 1270 285 1320 300
rect 1270 15 1285 285
rect 1305 15 1320 285
rect 1270 0 1320 15
rect 110 -120 160 -105
rect 110 -390 125 -120
rect 145 -390 160 -120
rect 110 -405 160 -390
rect 210 -120 260 -105
rect 210 -390 225 -120
rect 245 -390 260 -120
rect 210 -405 260 -390
rect 310 -120 360 -105
rect 310 -390 325 -120
rect 345 -390 360 -120
rect 310 -405 360 -390
rect 410 -120 460 -105
rect 410 -390 425 -120
rect 445 -390 460 -120
rect 410 -405 460 -390
rect 510 -120 560 -105
rect 510 -390 525 -120
rect 545 -390 560 -120
rect 510 -405 560 -390
rect 610 -120 660 -105
rect 610 -390 625 -120
rect 645 -390 660 -120
rect 610 -405 660 -390
rect 710 -120 760 -105
rect 710 -390 725 -120
rect 745 -390 760 -120
rect 710 -405 760 -390
rect 810 -120 860 -105
rect 810 -390 825 -120
rect 845 -390 860 -120
rect 810 -405 860 -390
rect 910 -120 960 -105
rect 910 -390 925 -120
rect 945 -390 960 -120
rect 910 -405 960 -390
rect 1010 -120 1060 -105
rect 1010 -390 1025 -120
rect 1045 -390 1060 -120
rect 1010 -405 1060 -390
rect 1110 -120 1160 -105
rect 1110 -390 1125 -120
rect 1145 -390 1160 -120
rect 1110 -405 1160 -390
<< pdiff >>
rect 110 1125 160 1140
rect 110 855 125 1125
rect 145 855 160 1125
rect 110 840 160 855
rect 210 1125 260 1140
rect 210 855 225 1125
rect 245 855 260 1125
rect 210 840 260 855
rect 310 1125 360 1140
rect 310 855 325 1125
rect 345 855 360 1125
rect 310 840 360 855
rect 410 1125 460 1140
rect 410 855 425 1125
rect 445 855 460 1125
rect 410 840 460 855
rect 510 1125 560 1140
rect 510 855 525 1125
rect 545 855 560 1125
rect 510 840 560 855
rect 610 1125 660 1140
rect 610 855 625 1125
rect 645 855 660 1125
rect 610 840 660 855
rect 710 1125 760 1140
rect 710 855 725 1125
rect 745 855 760 1125
rect 710 840 760 855
rect 810 1125 860 1140
rect 810 855 825 1125
rect 845 855 860 1125
rect 810 840 860 855
rect 910 1125 960 1140
rect 910 855 925 1125
rect 945 855 960 1125
rect 910 840 960 855
rect 1010 1125 1060 1140
rect 1010 855 1025 1125
rect 1045 855 1060 1125
rect 1010 840 1060 855
rect 1110 1125 1160 1140
rect 1110 855 1125 1125
rect 1145 855 1160 1125
rect 1110 840 1160 855
rect -50 680 0 695
rect -50 410 -35 680
rect -15 410 0 680
rect -50 395 0 410
rect 50 680 100 695
rect 50 410 65 680
rect 85 410 100 680
rect 50 395 100 410
rect 150 680 200 695
rect 150 410 165 680
rect 185 410 200 680
rect 150 395 200 410
rect 230 680 280 695
rect 230 410 245 680
rect 265 410 280 680
rect 230 395 280 410
rect 330 680 380 695
rect 330 410 345 680
rect 365 410 380 680
rect 330 395 380 410
rect 430 680 480 695
rect 430 410 445 680
rect 465 410 480 680
rect 430 395 480 410
rect 510 680 560 695
rect 510 410 525 680
rect 545 410 560 680
rect 510 395 560 410
rect 610 680 660 695
rect 610 410 625 680
rect 645 410 660 680
rect 610 395 660 410
rect 710 680 760 695
rect 710 410 725 680
rect 745 410 760 680
rect 710 395 760 410
rect 790 680 840 695
rect 790 410 805 680
rect 825 410 840 680
rect 790 395 840 410
rect 890 680 940 695
rect 890 410 905 680
rect 925 410 940 680
rect 890 395 940 410
rect 990 680 1040 695
rect 990 410 1005 680
rect 1025 410 1040 680
rect 990 395 1040 410
rect 1070 680 1120 695
rect 1070 410 1085 680
rect 1105 410 1120 680
rect 1070 395 1120 410
rect 1170 680 1220 695
rect 1170 410 1185 680
rect 1205 410 1220 680
rect 1170 395 1220 410
rect 1270 680 1320 695
rect 1270 410 1285 680
rect 1305 410 1320 680
rect 1270 395 1320 410
<< ndiffc >>
rect 125 1830 145 2100
rect 225 1830 245 2100
rect 325 1830 345 2100
rect 425 1830 445 2100
rect 525 1830 545 2100
rect 625 1830 645 2100
rect 725 1830 745 2100
rect 825 1830 845 2100
rect 925 1830 945 2100
rect 1025 1830 1045 2100
rect 1125 1830 1145 2100
rect 125 1360 145 1630
rect 225 1360 245 1630
rect 325 1360 345 1630
rect 425 1360 445 1630
rect 525 1360 545 1630
rect 625 1360 645 1630
rect 725 1360 745 1630
rect 825 1360 845 1630
rect 925 1360 945 1630
rect 1025 1360 1045 1630
rect 1125 1360 1145 1630
rect -35 15 -15 285
rect 65 15 85 285
rect 165 15 185 285
rect 245 15 265 285
rect 345 15 365 285
rect 445 15 465 285
rect 525 15 545 285
rect 625 15 645 285
rect 725 15 745 285
rect 805 15 825 285
rect 905 15 925 285
rect 1005 15 1025 285
rect 1085 15 1105 285
rect 1185 15 1205 285
rect 1285 15 1305 285
rect 125 -390 145 -120
rect 225 -390 245 -120
rect 325 -390 345 -120
rect 425 -390 445 -120
rect 525 -390 545 -120
rect 625 -390 645 -120
rect 725 -390 745 -120
rect 825 -390 845 -120
rect 925 -390 945 -120
rect 1025 -390 1045 -120
rect 1125 -390 1145 -120
<< pdiffc >>
rect 125 855 145 1125
rect 225 855 245 1125
rect 325 855 345 1125
rect 425 855 445 1125
rect 525 855 545 1125
rect 625 855 645 1125
rect 725 855 745 1125
rect 825 855 845 1125
rect 925 855 945 1125
rect 1025 855 1045 1125
rect 1125 855 1145 1125
rect -35 410 -15 680
rect 65 410 85 680
rect 165 410 185 680
rect 245 410 265 680
rect 345 410 365 680
rect 445 410 465 680
rect 525 410 545 680
rect 625 410 645 680
rect 725 410 745 680
rect 805 410 825 680
rect 905 410 925 680
rect 1005 410 1025 680
rect 1085 410 1105 680
rect 1185 410 1205 680
rect 1285 410 1305 680
<< poly >>
rect 160 2160 210 2170
rect 160 2140 175 2160
rect 195 2140 210 2160
rect 160 2115 210 2140
rect 260 2130 1010 2180
rect 260 2115 310 2130
rect 360 2115 410 2130
rect 460 2115 510 2130
rect 560 2115 610 2130
rect 660 2115 710 2130
rect 760 2115 810 2130
rect 860 2115 910 2130
rect 960 2115 1010 2130
rect 1060 2160 1110 2170
rect 1060 2140 1075 2160
rect 1095 2140 1110 2160
rect 1060 2115 1110 2140
rect 160 1800 210 1815
rect 260 1800 310 1815
rect 360 1800 410 1815
rect 460 1800 510 1815
rect 560 1800 610 1815
rect 660 1800 710 1815
rect 760 1800 810 1815
rect 860 1800 910 1815
rect 960 1800 1010 1815
rect 1060 1800 1110 1815
rect 110 1735 285 1775
rect 110 1725 910 1735
rect 160 1690 210 1700
rect 160 1670 175 1690
rect 195 1670 210 1690
rect 235 1685 910 1725
rect 160 1645 210 1670
rect 260 1645 310 1660
rect 360 1645 410 1685
rect 460 1645 510 1685
rect 560 1645 610 1660
rect 660 1645 710 1660
rect 760 1645 810 1685
rect 860 1645 910 1685
rect 1060 1690 1110 1700
rect 1060 1670 1075 1690
rect 1095 1670 1110 1690
rect 960 1645 1010 1660
rect 1060 1645 1110 1670
rect 160 1330 210 1345
rect 260 1305 310 1345
rect 360 1330 410 1345
rect 460 1330 510 1345
rect 560 1305 610 1345
rect 660 1305 710 1345
rect 760 1330 810 1345
rect 860 1330 910 1345
rect 960 1305 1010 1345
rect 1060 1330 1110 1345
rect 110 1255 1010 1305
rect 110 1205 310 1230
rect 110 1180 1010 1205
rect 260 1155 1010 1180
rect 160 1140 210 1155
rect 260 1140 310 1155
rect 360 1140 410 1155
rect 460 1140 510 1155
rect 560 1140 610 1155
rect 660 1140 710 1155
rect 760 1140 810 1155
rect 860 1140 910 1155
rect 960 1140 1010 1155
rect 1060 1140 1110 1155
rect -55 775 125 825
rect 160 815 210 840
rect 260 825 310 840
rect 360 825 410 840
rect 460 825 510 840
rect 560 825 610 840
rect 660 825 710 840
rect 760 825 810 840
rect 860 825 910 840
rect 960 825 1010 840
rect 160 795 175 815
rect 195 795 210 815
rect 160 785 210 795
rect 1060 815 1110 840
rect 1060 795 1075 815
rect 1095 795 1110 815
rect 1060 785 1110 795
rect 75 760 125 775
rect 0 740 50 750
rect 0 720 15 740
rect 35 720 50 740
rect 0 695 50 720
rect 75 710 1170 760
rect 100 695 150 710
rect 280 695 330 710
rect 380 695 430 710
rect 560 695 610 710
rect 660 695 710 710
rect 840 695 890 710
rect 940 695 990 710
rect 1120 695 1170 710
rect 1220 740 1270 750
rect 1220 720 1235 740
rect 1255 720 1270 740
rect 1220 695 1270 720
rect 0 380 50 395
rect 100 380 150 395
rect 280 380 330 395
rect 380 380 430 395
rect 560 380 610 395
rect 660 380 710 395
rect 840 380 890 395
rect 940 380 990 395
rect 1120 380 1170 395
rect 1220 380 1270 395
rect 475 345 805 355
rect 475 325 485 345
rect 505 340 775 345
rect 505 325 515 340
rect 475 315 515 325
rect 765 325 775 340
rect 795 325 805 345
rect 765 315 805 325
rect 0 300 50 315
rect 100 300 150 315
rect 280 300 330 315
rect 380 300 430 315
rect 560 300 610 315
rect 660 300 710 315
rect 840 300 890 315
rect 940 300 990 315
rect 1120 300 1170 315
rect 1220 300 1270 315
rect 0 -25 50 0
rect 0 -45 15 -25
rect 35 -45 50 -25
rect 0 -55 50 -45
rect 100 -15 150 0
rect 280 -15 330 0
rect 380 -15 430 0
rect 560 -15 610 0
rect 660 -15 710 0
rect 840 -15 890 0
rect 940 -15 990 0
rect 1120 -15 1170 0
rect 100 -65 1170 -15
rect 1220 -25 1270 0
rect 1220 -45 1235 -25
rect 1255 -45 1270 -25
rect 1220 -55 1270 -45
rect 160 -105 210 -90
rect 260 -105 310 -90
rect 360 -105 410 -90
rect 460 -105 510 -90
rect 560 -105 610 -90
rect 660 -105 710 -90
rect 760 -105 810 -90
rect 860 -105 910 -90
rect 960 -105 1010 -90
rect 1060 -105 1110 -90
rect 160 -430 210 -405
rect 160 -450 175 -430
rect 195 -450 210 -430
rect 160 -460 210 -450
rect 260 -420 310 -405
rect 360 -420 410 -405
rect 460 -420 510 -405
rect 560 -420 610 -405
rect 660 -420 710 -405
rect 760 -420 810 -405
rect 860 -420 910 -405
rect 960 -420 1010 -405
rect 260 -470 1010 -420
rect 1060 -430 1110 -405
rect 1060 -450 1075 -430
rect 1095 -450 1110 -430
rect 1060 -460 1110 -450
<< polycont >>
rect 175 2140 195 2160
rect 1075 2140 1095 2160
rect 175 1670 195 1690
rect 1075 1670 1095 1690
rect 175 795 195 815
rect 1075 795 1095 815
rect 15 720 35 740
rect 1235 720 1255 740
rect 485 325 505 345
rect 775 325 795 345
rect 15 -45 35 -25
rect 1235 -45 1255 -25
rect 175 -450 195 -430
rect 1075 -450 1095 -430
<< locali >>
rect 165 2160 205 2170
rect 165 2140 175 2160
rect 195 2140 205 2160
rect 165 2130 205 2140
rect 1065 2160 1105 2170
rect 1065 2140 1075 2160
rect 1095 2140 1105 2160
rect 1065 2130 1105 2140
rect 115 2100 155 2110
rect 115 1830 125 2100
rect 145 1830 155 2100
rect 115 1820 155 1830
rect 215 2100 255 2110
rect 215 1830 225 2100
rect 245 1830 255 2100
rect 215 1820 255 1830
rect 315 2100 355 2110
rect 315 1830 325 2100
rect 345 1830 355 2100
rect 315 1820 355 1830
rect 415 2100 455 2110
rect 415 1830 425 2100
rect 445 1830 455 2100
rect 415 1820 455 1830
rect 515 2100 555 2110
rect 515 1830 525 2100
rect 545 1830 555 2100
rect 515 1820 555 1830
rect 615 2100 655 2110
rect 615 1830 625 2100
rect 645 1830 655 2100
rect 615 1820 655 1830
rect 715 2100 755 2110
rect 715 1830 725 2100
rect 745 1830 755 2100
rect 715 1820 755 1830
rect 815 2100 855 2110
rect 815 1830 825 2100
rect 845 1830 855 2100
rect 815 1820 855 1830
rect 915 2100 955 2110
rect 915 1830 925 2100
rect 945 1830 955 2100
rect 915 1820 955 1830
rect 1015 2100 1055 2110
rect 1015 1830 1025 2100
rect 1045 1830 1055 2100
rect 1015 1820 1055 1830
rect 1115 2100 1155 2110
rect 1115 1830 1125 2100
rect 1145 1830 1155 2100
rect 1115 1820 1155 1830
rect 235 1740 255 1820
rect 425 1740 445 1820
rect 625 1740 645 1820
rect 825 1740 845 1820
rect 1015 1740 1035 1820
rect 235 1720 1035 1740
rect 165 1690 205 1700
rect 165 1670 175 1690
rect 195 1670 205 1690
rect 165 1660 205 1670
rect 325 1640 345 1720
rect 525 1640 545 1720
rect 725 1640 745 1720
rect 925 1640 945 1720
rect 1065 1690 1105 1700
rect 1065 1670 1075 1690
rect 1095 1670 1105 1690
rect 1065 1660 1105 1670
rect 115 1630 155 1640
rect 115 1360 125 1630
rect 145 1360 155 1630
rect 115 1350 155 1360
rect 215 1630 255 1640
rect 215 1360 225 1630
rect 245 1360 255 1630
rect 215 1350 255 1360
rect 315 1630 355 1640
rect 315 1360 325 1630
rect 345 1360 355 1630
rect 315 1350 355 1360
rect 415 1630 455 1640
rect 415 1360 425 1630
rect 445 1360 455 1630
rect 415 1350 455 1360
rect 515 1630 555 1640
rect 515 1360 525 1630
rect 545 1360 555 1630
rect 515 1350 555 1360
rect 615 1630 655 1640
rect 615 1360 625 1630
rect 645 1360 655 1630
rect 615 1350 655 1360
rect 715 1630 755 1640
rect 715 1360 725 1630
rect 745 1360 755 1630
rect 715 1350 755 1360
rect 815 1630 855 1640
rect 815 1360 825 1630
rect 845 1360 855 1630
rect 815 1350 855 1360
rect 915 1630 955 1640
rect 915 1360 925 1630
rect 945 1360 955 1630
rect 915 1350 955 1360
rect 1015 1630 1055 1640
rect 1015 1360 1025 1630
rect 1045 1360 1055 1630
rect 1015 1350 1055 1360
rect 1115 1630 1155 1640
rect 1115 1360 1125 1630
rect 1145 1360 1155 1630
rect 1115 1350 1155 1360
rect 225 1135 245 1350
rect 425 1135 445 1350
rect 625 1135 645 1350
rect 825 1135 845 1350
rect 1025 1135 1045 1350
rect 115 1125 155 1135
rect 115 855 125 1125
rect 145 855 155 1125
rect 115 845 155 855
rect 215 1125 255 1135
rect 215 855 225 1125
rect 245 855 255 1125
rect 215 845 255 855
rect 315 1125 355 1135
rect 315 855 325 1125
rect 345 855 355 1125
rect 315 845 355 855
rect 415 1125 455 1135
rect 415 855 425 1125
rect 445 855 455 1125
rect 415 845 455 855
rect 515 1125 555 1135
rect 515 855 525 1125
rect 545 855 555 1125
rect 515 845 555 855
rect 615 1125 655 1135
rect 615 855 625 1125
rect 645 855 655 1125
rect 615 845 655 855
rect 715 1125 755 1135
rect 715 855 725 1125
rect 745 855 755 1125
rect 715 845 755 855
rect 815 1125 855 1135
rect 815 855 825 1125
rect 845 855 855 1125
rect 815 845 855 855
rect 915 1125 955 1135
rect 915 855 925 1125
rect 945 855 955 1125
rect 915 845 955 855
rect 1015 1125 1055 1135
rect 1015 855 1025 1125
rect 1045 855 1055 1125
rect 1015 845 1055 855
rect 1115 1125 1155 1135
rect 1115 855 1125 1125
rect 1145 855 1155 1125
rect 1115 845 1155 855
rect 225 825 245 845
rect 425 825 445 845
rect 625 825 645 845
rect 825 825 845 845
rect 1025 825 1045 845
rect 165 815 205 825
rect 165 795 175 815
rect 195 795 205 815
rect 165 785 205 795
rect 1065 815 1105 825
rect 1065 795 1075 815
rect 1095 795 1105 815
rect 1065 785 1105 795
rect 5 740 45 750
rect 5 720 15 740
rect 35 720 45 740
rect 5 710 45 720
rect 1225 740 1265 750
rect 1225 720 1235 740
rect 1255 720 1265 740
rect 1225 710 1265 720
rect 65 690 85 710
rect 345 690 365 700
rect 625 690 645 700
rect 905 690 925 700
rect 1185 690 1205 700
rect -45 680 -5 690
rect -45 410 -35 680
rect -15 410 -5 680
rect -45 400 -5 410
rect 55 680 95 690
rect 55 410 65 680
rect 85 410 95 680
rect 55 400 95 410
rect 155 680 195 690
rect 155 410 165 680
rect 185 410 195 680
rect 155 400 195 410
rect 235 680 275 690
rect 235 410 245 680
rect 265 410 275 680
rect 235 400 275 410
rect 335 680 375 690
rect 335 410 345 680
rect 365 410 375 680
rect 335 400 375 410
rect 435 680 475 690
rect 435 410 445 680
rect 465 410 475 680
rect 435 400 475 410
rect 515 680 555 690
rect 515 410 525 680
rect 545 410 555 680
rect 515 400 555 410
rect 615 680 655 690
rect 615 410 625 680
rect 645 410 655 680
rect 615 400 655 410
rect 715 680 755 690
rect 715 410 725 680
rect 745 410 755 680
rect 715 400 755 410
rect 795 680 835 690
rect 795 410 805 680
rect 825 410 835 680
rect 795 400 835 410
rect 895 680 935 690
rect 895 410 905 680
rect 925 410 935 680
rect 895 400 935 410
rect 995 680 1035 690
rect 995 410 1005 680
rect 1025 410 1035 680
rect 995 400 1035 410
rect 1075 680 1115 690
rect 1075 410 1085 680
rect 1105 410 1115 680
rect 1075 400 1115 410
rect 1175 680 1215 690
rect 1175 410 1185 680
rect 1205 410 1215 680
rect 1175 400 1215 410
rect 1275 680 1315 690
rect 1275 410 1285 680
rect 1305 410 1315 680
rect 1275 400 1315 410
rect 175 355 195 400
rect 175 345 215 355
rect 175 325 185 345
rect 205 325 215 345
rect 175 315 215 325
rect 245 335 265 400
rect 455 355 475 400
rect 455 345 515 355
rect 455 335 485 345
rect 245 325 485 335
rect 505 325 515 345
rect 245 315 515 325
rect 535 335 555 400
rect 615 345 655 355
rect 615 335 625 345
rect 535 325 625 335
rect 645 335 655 345
rect 725 335 745 400
rect 805 355 825 400
rect 645 325 745 335
rect 535 315 745 325
rect 765 345 825 355
rect 765 325 775 345
rect 795 335 825 345
rect 1005 335 1025 400
rect 1075 355 1095 400
rect 795 325 1025 335
rect 765 315 1025 325
rect 1055 345 1095 355
rect 1055 325 1065 345
rect 1085 325 1095 345
rect 1055 315 1095 325
rect 175 295 195 315
rect 245 295 265 315
rect 455 295 475 315
rect 535 295 555 315
rect 725 295 745 315
rect 805 295 825 315
rect 1005 295 1025 315
rect 1075 295 1095 315
rect -45 285 -5 295
rect -45 15 -35 285
rect -15 15 -5 285
rect -45 5 -5 15
rect 55 285 95 295
rect 55 15 65 285
rect 85 15 95 285
rect 55 5 95 15
rect 155 285 195 295
rect 155 15 165 285
rect 185 15 195 285
rect 155 5 195 15
rect 235 285 275 295
rect 235 15 245 285
rect 265 15 275 285
rect 235 5 275 15
rect 335 285 375 295
rect 335 15 345 285
rect 365 15 375 285
rect 335 5 375 15
rect 435 285 475 295
rect 435 15 445 285
rect 465 15 475 285
rect 435 5 475 15
rect 515 285 555 295
rect 515 15 525 285
rect 545 15 555 285
rect 515 5 555 15
rect 615 285 655 295
rect 615 15 625 285
rect 645 15 655 285
rect 615 5 655 15
rect 715 285 755 295
rect 715 15 725 285
rect 745 15 755 285
rect 715 5 755 15
rect 795 285 835 295
rect 795 15 805 285
rect 825 15 835 285
rect 795 5 835 15
rect 895 285 935 295
rect 895 15 905 285
rect 925 15 935 285
rect 895 5 935 15
rect 995 285 1035 295
rect 995 15 1005 285
rect 1025 15 1035 285
rect 995 5 1035 15
rect 1075 285 1115 295
rect 1075 15 1085 285
rect 1105 15 1115 285
rect 1075 5 1115 15
rect 1175 285 1215 295
rect 1175 15 1185 285
rect 1205 15 1215 285
rect 1175 5 1215 15
rect 1275 285 1315 295
rect 1275 15 1285 285
rect 1305 15 1315 285
rect 1275 5 1315 15
rect 5 -25 45 -15
rect 5 -45 15 -25
rect 35 -45 45 -25
rect 5 -55 45 -45
rect 65 -70 85 5
rect 345 -70 365 5
rect 225 -110 245 -75
rect 425 -110 445 -70
rect 625 -110 645 5
rect 905 -75 925 5
rect 1185 -75 1205 5
rect 1225 -25 1265 -15
rect 1225 -45 1235 -25
rect 1255 -45 1265 -25
rect 1225 -55 1265 -45
rect 825 -110 845 -75
rect 1025 -110 1045 -75
rect 115 -120 155 -110
rect 115 -390 125 -120
rect 145 -390 155 -120
rect 115 -400 155 -390
rect 215 -120 255 -110
rect 215 -390 225 -120
rect 245 -390 255 -120
rect 215 -400 255 -390
rect 315 -120 355 -110
rect 315 -390 325 -120
rect 345 -390 355 -120
rect 315 -400 355 -390
rect 415 -120 455 -110
rect 415 -390 425 -120
rect 445 -390 455 -120
rect 415 -400 455 -390
rect 515 -120 555 -110
rect 515 -390 525 -120
rect 545 -390 555 -120
rect 515 -400 555 -390
rect 615 -120 655 -110
rect 615 -390 625 -120
rect 645 -390 655 -120
rect 615 -400 655 -390
rect 715 -120 755 -110
rect 715 -390 725 -120
rect 745 -390 755 -120
rect 715 -400 755 -390
rect 815 -120 855 -110
rect 815 -390 825 -120
rect 845 -390 855 -120
rect 815 -400 855 -390
rect 915 -120 955 -110
rect 915 -390 925 -120
rect 945 -390 955 -120
rect 915 -400 955 -390
rect 1015 -120 1055 -110
rect 1015 -390 1025 -120
rect 1045 -390 1055 -120
rect 1015 -400 1055 -390
rect 1115 -120 1155 -110
rect 1115 -390 1125 -120
rect 1145 -390 1155 -120
rect 1115 -400 1155 -390
rect 165 -430 205 -420
rect 165 -450 175 -430
rect 195 -450 205 -430
rect 165 -460 205 -450
rect 1065 -430 1105 -420
rect 1065 -450 1075 -430
rect 1095 -450 1105 -430
rect 1065 -460 1105 -450
<< viali >>
rect 125 1830 145 2100
rect 325 1830 345 2100
rect 525 1830 545 2100
rect 725 1830 745 2100
rect 925 1830 945 2100
rect 1125 1830 1145 2100
rect 125 1360 145 1630
rect 1125 1360 1145 1630
rect 125 855 145 1125
rect 325 855 345 1125
rect 525 855 545 1125
rect 725 855 745 1125
rect 925 855 945 1125
rect 1125 855 1145 1125
rect 185 325 205 345
rect 625 325 645 345
rect 1065 325 1085 345
rect 125 -390 145 -120
rect 325 -390 345 -120
rect 525 -390 545 -120
rect 725 -390 745 -120
rect 925 -390 945 -120
rect 1125 -390 1145 -120
<< metal1 >>
rect 175 345 1095 355
rect 175 325 185 345
rect 205 340 625 345
rect 205 325 215 340
rect 175 315 215 325
rect 615 325 625 340
rect 645 340 1065 345
rect 645 325 655 340
rect 615 315 655 325
rect 1055 325 1065 340
rect 1085 325 1095 345
rect 1055 315 1095 325
<< end >>
