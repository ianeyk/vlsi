** sch_path: /home/madvlsi/dev/git/vlsi/mp1/buffer/buffer.sch
**.subckt buffer VP VN A Y
*.iopin VP
*.iopin VN
*.ipin A
*.opin Y
x1 VP A net1 VN inverter
x2 VP net1 Y VN inverter
**.ends

* expanding   symbol:  /home/madvlsi/Documents/vlsi/mp1/inverter/inverter.sym # of pins=4
** sym_path: /home/madvlsi/Documents/vlsi/mp1/inverter/inverter.sym
** sch_path: /home/madvlsi/Documents/vlsi/mp1/inverter/inverter.sch
.subckt inverter VP A Y VN
*.iopin VP
*.iopin VN
*.ipin A
*.opin Y
XM1 Y A VN VN sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 Y A VP VP sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
