magic
tech sky130A
timestamp 1696998305
<< error_p >>
rect -35 2007 -15 2010
rect -35 1743 -32 2007
rect -18 1743 -15 2007
rect -35 1740 -15 1743
rect 165 2007 185 2010
rect 165 1743 168 2007
rect 182 1743 185 2007
rect 165 1740 185 1743
rect 245 2007 265 2010
rect 245 1743 248 2007
rect 262 1743 265 2007
rect 245 1740 265 1743
rect 445 2007 465 2010
rect 445 1743 448 2007
rect 462 1743 465 2007
rect 445 1740 465 1743
rect 525 2007 545 2010
rect 525 1743 528 2007
rect 542 1743 545 2007
rect 525 1740 545 1743
rect 725 2007 745 2010
rect 725 1743 728 2007
rect 742 1743 745 2007
rect 725 1740 745 1743
rect 805 2007 825 2010
rect 805 1743 808 2007
rect 822 1743 825 2007
rect 805 1740 825 1743
rect 1005 2007 1025 2010
rect 1005 1743 1008 2007
rect 1022 1743 1025 2007
rect 1005 1740 1025 1743
rect 1085 2007 1105 2010
rect 1085 1743 1088 2007
rect 1102 1743 1105 2007
rect 1085 1740 1105 1743
rect 1285 2007 1305 2010
rect 1285 1743 1288 2007
rect 1302 1743 1305 2007
rect 1285 1740 1305 1743
rect -35 1537 -15 1540
rect -35 1273 -32 1537
rect -18 1273 -15 1537
rect -35 1270 -15 1273
rect 1285 1537 1305 1540
rect 1285 1273 1288 1537
rect 1302 1273 1305 1537
rect 1285 1270 1305 1273
rect -35 1057 -15 1060
rect -35 793 -32 1057
rect -18 793 -15 1057
rect -35 790 -15 793
rect 165 1057 185 1060
rect 165 793 168 1057
rect 182 793 185 1057
rect 165 790 185 793
rect 245 1057 265 1060
rect 245 793 248 1057
rect 262 793 265 1057
rect 245 790 265 793
rect 445 1057 465 1060
rect 445 793 448 1057
rect 462 793 465 1057
rect 445 790 465 793
rect 525 1057 545 1060
rect 525 793 528 1057
rect 542 793 545 1057
rect 525 790 545 793
rect 725 1057 745 1060
rect 725 793 728 1057
rect 742 793 745 1057
rect 725 790 745 793
rect 805 1057 825 1060
rect 805 793 808 1057
rect 822 793 825 1057
rect 805 790 825 793
rect 1005 1057 1025 1060
rect 1005 793 1008 1057
rect 1022 793 1025 1057
rect 1005 790 1025 793
rect 1085 1057 1105 1060
rect 1085 793 1088 1057
rect 1102 793 1105 1057
rect 1085 790 1105 793
rect 1285 1057 1305 1060
rect 1285 793 1288 1057
rect 1302 793 1305 1057
rect 1285 790 1305 793
rect -35 -123 -15 -120
rect -35 -387 -32 -123
rect -18 -387 -15 -123
rect -35 -390 -15 -387
rect 165 -123 185 -120
rect 165 -387 168 -123
rect 182 -387 185 -123
rect 165 -390 185 -387
rect 245 -123 265 -120
rect 245 -387 248 -123
rect 262 -387 265 -123
rect 245 -390 265 -387
rect 445 -123 465 -120
rect 445 -387 448 -123
rect 462 -387 465 -123
rect 445 -390 465 -387
rect 525 -123 545 -120
rect 525 -387 528 -123
rect 542 -387 545 -123
rect 525 -390 545 -387
rect 725 -123 745 -120
rect 725 -387 728 -123
rect 742 -387 745 -123
rect 725 -390 745 -387
rect 805 -123 825 -120
rect 805 -387 808 -123
rect 822 -387 825 -123
rect 805 -390 825 -387
rect 1005 -123 1025 -120
rect 1005 -387 1008 -123
rect 1022 -387 1025 -123
rect 1005 -390 1025 -387
rect 1085 -123 1105 -120
rect 1085 -387 1088 -123
rect 1102 -387 1105 -123
rect 1085 -390 1105 -387
rect 1285 -123 1305 -120
rect 1285 -387 1288 -123
rect 1302 -387 1305 -123
rect 1285 -390 1305 -387
<< nwell >>
rect -70 335 1340 1095
<< nmos >>
rect 0 1725 50 2025
rect 100 1725 150 2025
rect 280 1725 330 2025
rect 380 1725 430 2025
rect 560 1725 610 2025
rect 660 1725 710 2025
rect 840 1725 890 2025
rect 940 1725 990 2025
rect 1120 1725 1170 2025
rect 1220 1725 1270 2025
rect 0 1255 50 1555
rect 100 1255 150 1555
rect 280 1255 330 1555
rect 380 1255 430 1555
rect 560 1255 610 1555
rect 660 1255 710 1555
rect 840 1255 890 1555
rect 940 1255 990 1555
rect 1120 1255 1170 1555
rect 1220 1255 1270 1555
rect 0 0 50 300
rect 100 0 150 300
rect 280 0 330 300
rect 380 0 430 300
rect 560 0 610 300
rect 660 0 710 300
rect 840 0 890 300
rect 940 0 990 300
rect 1120 0 1170 300
rect 1220 0 1270 300
rect 0 -405 50 -105
rect 100 -405 150 -105
rect 280 -405 330 -105
rect 380 -405 430 -105
rect 560 -405 610 -105
rect 660 -405 710 -105
rect 840 -405 890 -105
rect 940 -405 990 -105
rect 1120 -405 1170 -105
rect 1220 -405 1270 -105
<< pmos >>
rect 0 775 50 1075
rect 100 775 150 1075
rect 280 775 330 1075
rect 380 775 430 1075
rect 560 775 610 1075
rect 660 775 710 1075
rect 840 775 890 1075
rect 940 775 990 1075
rect 1120 775 1170 1075
rect 1220 775 1270 1075
rect 0 355 50 655
rect 100 355 150 655
rect 280 355 330 655
rect 380 355 430 655
rect 560 355 610 655
rect 660 355 710 655
rect 840 355 890 655
rect 940 355 990 655
rect 1120 355 1170 655
rect 1220 355 1270 655
<< ndiff >>
rect -50 2010 0 2025
rect -50 1740 -35 2010
rect -15 1740 0 2010
rect -50 1725 0 1740
rect 50 2010 100 2025
rect 50 1740 65 2010
rect 85 1740 100 2010
rect 50 1725 100 1740
rect 150 2010 200 2025
rect 150 1740 165 2010
rect 185 1740 200 2010
rect 150 1725 200 1740
rect 230 2010 280 2025
rect 230 1740 245 2010
rect 265 1740 280 2010
rect 230 1725 280 1740
rect 330 2010 380 2025
rect 330 1740 345 2010
rect 365 1740 380 2010
rect 330 1725 380 1740
rect 430 2010 480 2025
rect 430 1740 445 2010
rect 465 1740 480 2010
rect 430 1725 480 1740
rect 510 2010 560 2025
rect 510 1740 525 2010
rect 545 1740 560 2010
rect 510 1725 560 1740
rect 610 2010 660 2025
rect 610 1740 625 2010
rect 645 1740 660 2010
rect 610 1725 660 1740
rect 710 2010 760 2025
rect 710 1740 725 2010
rect 745 1740 760 2010
rect 710 1725 760 1740
rect 790 2010 840 2025
rect 790 1740 805 2010
rect 825 1740 840 2010
rect 790 1725 840 1740
rect 890 2010 940 2025
rect 890 1740 905 2010
rect 925 1740 940 2010
rect 890 1725 940 1740
rect 990 2010 1040 2025
rect 990 1740 1005 2010
rect 1025 1740 1040 2010
rect 990 1725 1040 1740
rect 1070 2010 1120 2025
rect 1070 1740 1085 2010
rect 1105 1740 1120 2010
rect 1070 1725 1120 1740
rect 1170 2010 1220 2025
rect 1170 1740 1185 2010
rect 1205 1740 1220 2010
rect 1170 1725 1220 1740
rect 1270 2010 1320 2025
rect 1270 1740 1285 2010
rect 1305 1740 1320 2010
rect 1270 1725 1320 1740
rect -50 1540 0 1555
rect -50 1270 -35 1540
rect -15 1270 0 1540
rect -50 1255 0 1270
rect 50 1540 100 1555
rect 50 1270 65 1540
rect 85 1270 100 1540
rect 50 1255 100 1270
rect 150 1540 200 1555
rect 150 1270 165 1540
rect 185 1270 200 1540
rect 150 1255 200 1270
rect 230 1540 280 1555
rect 230 1270 245 1540
rect 265 1270 280 1540
rect 230 1255 280 1270
rect 330 1540 380 1555
rect 330 1270 345 1540
rect 365 1270 380 1540
rect 330 1255 380 1270
rect 430 1540 480 1555
rect 430 1270 445 1540
rect 465 1270 480 1540
rect 430 1255 480 1270
rect 510 1540 560 1555
rect 510 1270 525 1540
rect 545 1270 560 1540
rect 510 1255 560 1270
rect 610 1540 660 1555
rect 610 1270 625 1540
rect 645 1270 660 1540
rect 610 1255 660 1270
rect 710 1540 760 1555
rect 710 1270 725 1540
rect 745 1270 760 1540
rect 710 1255 760 1270
rect 790 1540 840 1555
rect 790 1270 805 1540
rect 825 1270 840 1540
rect 790 1255 840 1270
rect 890 1540 940 1555
rect 890 1270 905 1540
rect 925 1270 940 1540
rect 890 1255 940 1270
rect 990 1540 1040 1555
rect 990 1270 1005 1540
rect 1025 1270 1040 1540
rect 990 1255 1040 1270
rect 1070 1540 1120 1555
rect 1070 1270 1085 1540
rect 1105 1270 1120 1540
rect 1070 1255 1120 1270
rect 1170 1540 1220 1555
rect 1170 1270 1185 1540
rect 1205 1270 1220 1540
rect 1170 1255 1220 1270
rect 1270 1540 1320 1555
rect 1270 1270 1285 1540
rect 1305 1270 1320 1540
rect 1270 1255 1320 1270
rect -50 285 0 300
rect -50 15 -35 285
rect -15 15 0 285
rect -50 0 0 15
rect 50 285 100 300
rect 50 15 65 285
rect 85 15 100 285
rect 50 0 100 15
rect 150 285 200 300
rect 150 15 165 285
rect 185 15 200 285
rect 150 0 200 15
rect 230 285 280 300
rect 230 15 245 285
rect 265 15 280 285
rect 230 0 280 15
rect 330 285 380 300
rect 330 15 345 285
rect 365 15 380 285
rect 330 0 380 15
rect 430 285 480 300
rect 430 15 445 285
rect 465 15 480 285
rect 430 0 480 15
rect 510 285 560 300
rect 510 15 525 285
rect 545 15 560 285
rect 510 0 560 15
rect 610 285 660 300
rect 610 15 625 285
rect 645 15 660 285
rect 610 0 660 15
rect 710 285 760 300
rect 710 15 725 285
rect 745 15 760 285
rect 710 0 760 15
rect 790 285 840 300
rect 790 15 805 285
rect 825 15 840 285
rect 790 0 840 15
rect 890 285 940 300
rect 890 15 905 285
rect 925 15 940 285
rect 890 0 940 15
rect 990 285 1040 300
rect 990 15 1005 285
rect 1025 15 1040 285
rect 990 0 1040 15
rect 1070 285 1120 300
rect 1070 15 1085 285
rect 1105 15 1120 285
rect 1070 0 1120 15
rect 1170 285 1220 300
rect 1170 15 1185 285
rect 1205 15 1220 285
rect 1170 0 1220 15
rect 1270 285 1320 300
rect 1270 15 1285 285
rect 1305 15 1320 285
rect 1270 0 1320 15
rect -50 -120 0 -105
rect -50 -390 -35 -120
rect -15 -390 0 -120
rect -50 -405 0 -390
rect 50 -120 100 -105
rect 50 -390 65 -120
rect 85 -390 100 -120
rect 50 -405 100 -390
rect 150 -120 200 -105
rect 150 -390 165 -120
rect 185 -390 200 -120
rect 150 -405 200 -390
rect 230 -120 280 -105
rect 230 -390 245 -120
rect 265 -390 280 -120
rect 230 -405 280 -390
rect 330 -120 380 -105
rect 330 -390 345 -120
rect 365 -390 380 -120
rect 330 -405 380 -390
rect 430 -120 480 -105
rect 430 -390 445 -120
rect 465 -390 480 -120
rect 430 -405 480 -390
rect 510 -120 560 -105
rect 510 -390 525 -120
rect 545 -390 560 -120
rect 510 -405 560 -390
rect 610 -120 660 -105
rect 610 -390 625 -120
rect 645 -390 660 -120
rect 610 -405 660 -390
rect 710 -120 760 -105
rect 710 -390 725 -120
rect 745 -390 760 -120
rect 710 -405 760 -390
rect 790 -120 840 -105
rect 790 -390 805 -120
rect 825 -390 840 -120
rect 790 -405 840 -390
rect 890 -120 940 -105
rect 890 -390 905 -120
rect 925 -390 940 -120
rect 890 -405 940 -390
rect 990 -120 1040 -105
rect 990 -390 1005 -120
rect 1025 -390 1040 -120
rect 990 -405 1040 -390
rect 1070 -120 1120 -105
rect 1070 -390 1085 -120
rect 1105 -390 1120 -120
rect 1070 -405 1120 -390
rect 1170 -120 1220 -105
rect 1170 -390 1185 -120
rect 1205 -390 1220 -120
rect 1170 -405 1220 -390
rect 1270 -120 1320 -105
rect 1270 -390 1285 -120
rect 1305 -390 1320 -120
rect 1270 -405 1320 -390
<< pdiff >>
rect -50 1060 0 1075
rect -50 790 -35 1060
rect -15 790 0 1060
rect -50 775 0 790
rect 50 1060 100 1075
rect 50 790 65 1060
rect 85 790 100 1060
rect 50 775 100 790
rect 150 1060 200 1075
rect 150 790 165 1060
rect 185 790 200 1060
rect 150 775 200 790
rect 230 1060 280 1075
rect 230 790 245 1060
rect 265 790 280 1060
rect 230 775 280 790
rect 330 1060 380 1075
rect 330 790 345 1060
rect 365 790 380 1060
rect 330 775 380 790
rect 430 1060 480 1075
rect 430 790 445 1060
rect 465 790 480 1060
rect 430 775 480 790
rect 510 1060 560 1075
rect 510 790 525 1060
rect 545 790 560 1060
rect 510 775 560 790
rect 610 1060 660 1075
rect 610 790 625 1060
rect 645 790 660 1060
rect 610 775 660 790
rect 710 1060 760 1075
rect 710 790 725 1060
rect 745 790 760 1060
rect 710 775 760 790
rect 790 1060 840 1075
rect 790 790 805 1060
rect 825 790 840 1060
rect 790 775 840 790
rect 890 1060 940 1075
rect 890 790 905 1060
rect 925 790 940 1060
rect 890 775 940 790
rect 990 1060 1040 1075
rect 990 790 1005 1060
rect 1025 790 1040 1060
rect 990 775 1040 790
rect 1070 1060 1120 1075
rect 1070 790 1085 1060
rect 1105 790 1120 1060
rect 1070 775 1120 790
rect 1170 1060 1220 1075
rect 1170 790 1185 1060
rect 1205 790 1220 1060
rect 1170 775 1220 790
rect 1270 1060 1320 1075
rect 1270 790 1285 1060
rect 1305 790 1320 1060
rect 1270 775 1320 790
rect -50 640 0 655
rect -50 370 -35 640
rect -15 370 0 640
rect -50 355 0 370
rect 50 640 100 655
rect 50 370 65 640
rect 85 370 100 640
rect 50 355 100 370
rect 150 640 200 655
rect 150 370 165 640
rect 185 370 200 640
rect 150 355 200 370
rect 230 640 280 655
rect 230 370 245 640
rect 265 370 280 640
rect 230 355 280 370
rect 330 640 380 655
rect 330 370 345 640
rect 365 370 380 640
rect 330 355 380 370
rect 430 640 480 655
rect 430 370 445 640
rect 465 370 480 640
rect 430 355 480 370
rect 510 640 560 655
rect 510 370 525 640
rect 545 370 560 640
rect 510 355 560 370
rect 610 640 660 655
rect 610 370 625 640
rect 645 370 660 640
rect 610 355 660 370
rect 710 640 760 655
rect 710 370 725 640
rect 745 370 760 640
rect 710 355 760 370
rect 790 640 840 655
rect 790 370 805 640
rect 825 370 840 640
rect 790 355 840 370
rect 890 640 940 655
rect 890 370 905 640
rect 925 370 940 640
rect 890 355 940 370
rect 990 640 1040 655
rect 990 370 1005 640
rect 1025 370 1040 640
rect 990 355 1040 370
rect 1070 640 1120 655
rect 1070 370 1085 640
rect 1105 370 1120 640
rect 1070 355 1120 370
rect 1170 640 1220 655
rect 1170 370 1185 640
rect 1205 370 1220 640
rect 1170 355 1220 370
rect 1270 640 1320 655
rect 1270 370 1285 640
rect 1305 370 1320 640
rect 1270 355 1320 370
<< ndiffc >>
rect -35 1740 -15 2010
rect 65 1740 85 2010
rect 165 1740 185 2010
rect 245 1740 265 2010
rect 345 1740 365 2010
rect 445 1740 465 2010
rect 525 1740 545 2010
rect 625 1740 645 2010
rect 725 1740 745 2010
rect 805 1740 825 2010
rect 905 1740 925 2010
rect 1005 1740 1025 2010
rect 1085 1740 1105 2010
rect 1185 1740 1205 2010
rect 1285 1740 1305 2010
rect -35 1270 -15 1540
rect 65 1270 85 1540
rect 165 1270 185 1540
rect 245 1270 265 1540
rect 345 1270 365 1540
rect 445 1270 465 1540
rect 525 1270 545 1540
rect 625 1270 645 1540
rect 725 1270 745 1540
rect 805 1270 825 1540
rect 905 1270 925 1540
rect 1005 1270 1025 1540
rect 1085 1270 1105 1540
rect 1185 1270 1205 1540
rect 1285 1270 1305 1540
rect -35 15 -15 285
rect 65 15 85 285
rect 165 15 185 285
rect 245 15 265 285
rect 345 15 365 285
rect 445 15 465 285
rect 525 15 545 285
rect 625 15 645 285
rect 725 15 745 285
rect 805 15 825 285
rect 905 15 925 285
rect 1005 15 1025 285
rect 1085 15 1105 285
rect 1185 15 1205 285
rect 1285 15 1305 285
rect -35 -390 -15 -120
rect 65 -390 85 -120
rect 165 -390 185 -120
rect 245 -390 265 -120
rect 345 -390 365 -120
rect 445 -390 465 -120
rect 525 -390 545 -120
rect 625 -390 645 -120
rect 725 -390 745 -120
rect 805 -390 825 -120
rect 905 -390 925 -120
rect 1005 -390 1025 -120
rect 1085 -390 1105 -120
rect 1185 -390 1205 -120
rect 1285 -390 1305 -120
<< pdiffc >>
rect -35 790 -15 1060
rect 65 790 85 1060
rect 165 790 185 1060
rect 245 790 265 1060
rect 345 790 365 1060
rect 445 790 465 1060
rect 525 790 545 1060
rect 625 790 645 1060
rect 725 790 745 1060
rect 805 790 825 1060
rect 905 790 925 1060
rect 1005 790 1025 1060
rect 1085 790 1105 1060
rect 1185 790 1205 1060
rect 1285 790 1305 1060
rect -35 370 -15 640
rect 65 370 85 640
rect 165 370 185 640
rect 245 370 265 640
rect 345 370 365 640
rect 445 370 465 640
rect 525 370 545 640
rect 625 370 645 640
rect 725 370 745 640
rect 805 370 825 640
rect 905 370 925 640
rect 1005 370 1025 640
rect 1085 370 1105 640
rect 1185 370 1205 640
rect 1285 370 1305 640
<< poly >>
rect 0 2070 50 2080
rect 0 2050 15 2070
rect 35 2050 50 2070
rect 0 2025 50 2050
rect 100 2040 1170 2090
rect 100 2025 150 2040
rect 280 2025 330 2040
rect 380 2025 430 2040
rect 560 2025 610 2040
rect 660 2025 710 2040
rect 840 2025 890 2040
rect 940 2025 990 2040
rect 1120 2025 1170 2040
rect 1220 2070 1270 2080
rect 1220 2050 1235 2070
rect 1255 2050 1270 2070
rect 1220 2025 1270 2050
rect 0 1710 50 1725
rect 100 1710 150 1725
rect 280 1710 330 1725
rect 380 1710 430 1725
rect 560 1710 610 1725
rect 660 1710 710 1725
rect 840 1710 890 1725
rect 940 1710 990 1725
rect 1120 1710 1170 1725
rect 1220 1710 1270 1725
rect -50 1645 125 1685
rect -50 1635 990 1645
rect 0 1600 50 1610
rect 0 1580 15 1600
rect 35 1580 50 1600
rect 75 1595 990 1635
rect 0 1555 50 1580
rect 100 1555 150 1570
rect 280 1555 330 1595
rect 380 1555 430 1595
rect 560 1555 610 1570
rect 660 1555 710 1570
rect 840 1555 890 1595
rect 940 1555 990 1595
rect 1120 1555 1170 1570
rect 1220 1555 1270 1570
rect 0 1240 50 1255
rect 100 1215 150 1255
rect 280 1240 330 1255
rect 380 1240 430 1255
rect 560 1215 610 1255
rect 660 1215 710 1255
rect 840 1240 890 1255
rect 940 1240 990 1255
rect 1120 1215 1170 1255
rect -50 1165 1170 1215
rect 1220 1230 1270 1255
rect 1220 1210 1235 1230
rect 1255 1210 1270 1230
rect 1220 1200 1270 1210
rect 0 1120 50 1130
rect 0 1100 15 1120
rect 35 1100 50 1120
rect 0 1075 50 1100
rect 100 1090 1170 1140
rect 100 1075 150 1090
rect 280 1075 330 1090
rect 380 1075 430 1090
rect 560 1075 610 1090
rect 660 1075 710 1090
rect 840 1075 890 1090
rect 940 1075 990 1090
rect 1120 1075 1170 1090
rect 1220 1120 1270 1130
rect 1220 1100 1235 1120
rect 1255 1100 1270 1120
rect 1220 1075 1270 1100
rect 0 760 50 775
rect 100 760 150 775
rect 280 760 330 775
rect 380 760 430 775
rect 560 760 610 775
rect 660 760 710 775
rect 840 760 890 775
rect 940 760 990 775
rect 1120 760 1170 775
rect 1220 760 1270 775
rect 0 700 50 710
rect 0 680 15 700
rect 35 680 50 700
rect 0 655 50 680
rect 100 670 1170 720
rect 100 655 150 670
rect 280 655 330 670
rect 380 655 430 670
rect 560 655 610 670
rect 660 655 710 670
rect 840 655 890 670
rect 940 655 990 670
rect 1120 655 1170 670
rect 1220 700 1270 710
rect 1220 680 1235 700
rect 1255 680 1270 700
rect 1220 655 1270 680
rect 0 340 50 355
rect 100 340 150 355
rect 280 340 330 355
rect 380 340 430 355
rect 560 340 610 355
rect 660 340 710 355
rect 840 340 890 355
rect 940 340 990 355
rect 1120 340 1170 355
rect 1220 340 1270 355
rect 0 300 50 315
rect 100 300 150 315
rect 280 300 330 315
rect 380 300 430 315
rect 560 300 610 315
rect 660 300 710 315
rect 840 300 890 315
rect 940 300 990 315
rect 1120 300 1170 315
rect 1220 300 1270 315
rect 0 -25 50 0
rect 0 -45 15 -25
rect 35 -45 50 -25
rect 0 -55 50 -45
rect 100 -15 150 0
rect 280 -15 330 0
rect 380 -15 430 0
rect 560 -15 610 0
rect 660 -15 710 0
rect 840 -15 890 0
rect 940 -15 990 0
rect 1120 -15 1170 0
rect 100 -65 1170 -15
rect 1220 -25 1270 0
rect 1220 -45 1235 -25
rect 1255 -45 1270 -25
rect 1220 -55 1270 -45
rect 0 -105 50 -90
rect 100 -105 150 -90
rect 280 -105 330 -90
rect 380 -105 430 -90
rect 560 -105 610 -90
rect 660 -105 710 -90
rect 840 -105 890 -90
rect 940 -105 990 -90
rect 1120 -105 1170 -90
rect 1220 -105 1270 -90
rect 0 -430 50 -405
rect 0 -450 15 -430
rect 35 -450 50 -430
rect 0 -460 50 -450
rect 100 -420 150 -405
rect 280 -420 330 -405
rect 380 -420 430 -405
rect 560 -420 610 -405
rect 660 -420 710 -405
rect 840 -420 890 -405
rect 940 -420 990 -405
rect 1120 -420 1170 -405
rect 100 -470 1170 -420
rect 1220 -430 1270 -405
rect 1220 -450 1235 -430
rect 1255 -450 1270 -430
rect 1220 -460 1270 -450
<< polycont >>
rect 15 2050 35 2070
rect 1235 2050 1255 2070
rect 15 1580 35 1600
rect 1235 1210 1255 1230
rect 15 1100 35 1120
rect 1235 1100 1255 1120
rect 15 680 35 700
rect 1235 680 1255 700
rect 15 -45 35 -25
rect 1235 -45 1255 -25
rect 15 -450 35 -430
rect 1235 -450 1255 -430
<< locali >>
rect 5 2070 45 2080
rect 5 2050 15 2070
rect 35 2050 45 2070
rect 5 2040 45 2050
rect 1225 2070 1265 2080
rect 1225 2050 1235 2070
rect 1255 2050 1265 2070
rect 1225 2040 1265 2050
rect -45 2010 -5 2020
rect -45 1740 -35 2010
rect -15 1740 -5 2010
rect -45 1730 -5 1740
rect 55 2010 95 2020
rect 55 1740 65 2010
rect 85 1740 95 2010
rect 55 1730 95 1740
rect 155 2010 275 2020
rect 155 1740 165 2010
rect 185 1740 245 2010
rect 265 1740 275 2010
rect 155 1730 275 1740
rect 335 2010 375 2020
rect 335 1740 345 2010
rect 365 1740 375 2010
rect 335 1730 375 1740
rect 435 2010 555 2020
rect 435 1740 445 2010
rect 465 1740 525 2010
rect 545 1740 555 2010
rect 435 1730 555 1740
rect 615 2010 655 2020
rect 615 1740 625 2010
rect 645 1740 655 2010
rect 615 1730 655 1740
rect 715 2010 835 2020
rect 715 1740 725 2010
rect 745 1740 805 2010
rect 825 1740 835 2010
rect 715 1730 835 1740
rect 895 2010 935 2020
rect 895 1740 905 2010
rect 925 1740 935 2010
rect 895 1730 935 1740
rect 995 2010 1115 2020
rect 995 1740 1005 2010
rect 1025 1740 1085 2010
rect 1105 1740 1115 2010
rect 995 1730 1115 1740
rect 1175 2010 1215 2020
rect 1175 1740 1185 2010
rect 1205 1740 1215 2010
rect 1175 1730 1215 1740
rect 1275 2010 1315 2020
rect 1275 1740 1285 2010
rect 1305 1740 1315 2010
rect 1275 1730 1315 1740
rect 5 1600 45 1610
rect 5 1580 15 1600
rect 35 1580 45 1600
rect 5 1570 45 1580
rect -45 1540 -5 1550
rect -45 1270 -35 1540
rect -15 1270 -5 1540
rect -45 1260 -5 1270
rect 55 1540 95 1550
rect 55 1270 65 1540
rect 85 1270 95 1540
rect 55 1260 95 1270
rect 155 1540 195 1550
rect 155 1270 165 1540
rect 185 1270 195 1540
rect 155 1260 195 1270
rect 235 1540 275 1550
rect 235 1270 245 1540
rect 265 1270 275 1540
rect 235 1260 275 1270
rect 335 1540 375 1550
rect 335 1270 345 1540
rect 365 1270 375 1540
rect 335 1260 375 1270
rect 435 1540 475 1550
rect 435 1270 445 1540
rect 465 1270 475 1540
rect 435 1260 475 1270
rect 515 1540 555 1550
rect 515 1270 525 1540
rect 545 1270 555 1540
rect 515 1260 555 1270
rect 615 1540 655 1550
rect 615 1270 625 1540
rect 645 1270 655 1540
rect 615 1260 655 1270
rect 715 1540 755 1550
rect 715 1270 725 1540
rect 745 1270 755 1540
rect 715 1260 755 1270
rect 795 1540 835 1550
rect 795 1270 805 1540
rect 825 1270 835 1540
rect 795 1260 835 1270
rect 895 1540 935 1550
rect 895 1270 905 1540
rect 925 1270 935 1540
rect 895 1260 935 1270
rect 995 1540 1035 1550
rect 995 1270 1005 1540
rect 1025 1270 1035 1540
rect 995 1260 1035 1270
rect 1075 1540 1115 1550
rect 1075 1270 1085 1540
rect 1105 1270 1115 1540
rect 1075 1260 1115 1270
rect 1175 1540 1215 1550
rect 1175 1270 1185 1540
rect 1205 1270 1215 1540
rect 1175 1260 1215 1270
rect 1275 1540 1315 1550
rect 1275 1270 1285 1540
rect 1305 1270 1315 1540
rect 1275 1260 1315 1270
rect 65 1230 85 1260
rect 345 1230 365 1260
rect 625 1230 645 1260
rect 905 1230 925 1260
rect 1185 1230 1205 1260
rect 1225 1230 1265 1240
rect 1225 1210 1235 1230
rect 1255 1210 1265 1230
rect 1225 1200 1265 1210
rect 5 1120 45 1130
rect 5 1100 15 1120
rect 35 1100 45 1120
rect 1225 1120 1265 1130
rect 5 1090 45 1100
rect 65 1070 85 1105
rect 345 1070 365 1105
rect 625 1070 645 1105
rect 905 1070 925 1105
rect 1185 1070 1205 1105
rect 1225 1100 1235 1120
rect 1255 1100 1265 1120
rect 1225 1090 1265 1100
rect -45 1060 -5 1070
rect -45 790 -35 1060
rect -15 790 -5 1060
rect -45 780 -5 790
rect 55 1060 95 1070
rect 55 790 65 1060
rect 85 790 95 1060
rect 55 780 95 790
rect 155 1060 275 1070
rect 155 790 165 1060
rect 185 790 245 1060
rect 265 790 275 1060
rect 155 780 275 790
rect 335 1060 375 1070
rect 335 790 345 1060
rect 365 790 375 1060
rect 335 780 375 790
rect 435 1060 555 1070
rect 435 790 445 1060
rect 465 790 525 1060
rect 545 790 555 1060
rect 435 780 555 790
rect 615 1060 655 1070
rect 615 790 625 1060
rect 645 790 655 1060
rect 615 780 655 790
rect 715 1060 835 1070
rect 715 790 725 1060
rect 745 790 805 1060
rect 825 790 835 1060
rect 715 780 835 790
rect 895 1060 935 1070
rect 895 790 905 1060
rect 925 790 935 1060
rect 895 780 935 790
rect 995 1060 1115 1070
rect 995 790 1005 1060
rect 1025 790 1085 1060
rect 1105 790 1115 1060
rect 995 780 1115 790
rect 1175 1060 1215 1070
rect 1175 790 1185 1060
rect 1205 790 1215 1060
rect 1175 780 1215 790
rect 1275 1060 1315 1070
rect 1275 790 1285 1060
rect 1305 790 1315 1060
rect 1275 780 1315 790
rect 65 760 85 780
rect 345 760 365 780
rect 625 760 645 780
rect 905 760 925 780
rect 1185 760 1205 780
rect 5 700 45 710
rect 5 680 15 700
rect 35 680 45 700
rect 5 670 45 680
rect 1225 700 1265 710
rect 1225 680 1235 700
rect 1255 680 1265 700
rect 1225 670 1265 680
rect 65 650 85 670
rect 345 650 365 660
rect 625 650 645 660
rect 905 650 925 660
rect 1185 650 1205 660
rect -45 640 -5 650
rect -45 370 -35 640
rect -15 370 -5 640
rect -45 360 -5 370
rect 55 640 95 650
rect 55 370 65 640
rect 85 370 95 640
rect 55 360 95 370
rect 155 640 195 650
rect 155 370 165 640
rect 185 370 195 640
rect 155 360 195 370
rect 235 640 275 650
rect 235 370 245 640
rect 265 370 275 640
rect 235 360 275 370
rect 335 640 375 650
rect 335 370 345 640
rect 365 370 375 640
rect 335 360 375 370
rect 435 640 475 650
rect 435 370 445 640
rect 465 370 475 640
rect 435 360 475 370
rect 515 640 555 650
rect 515 370 525 640
rect 545 370 555 640
rect 515 360 555 370
rect 615 640 655 650
rect 615 370 625 640
rect 645 370 655 640
rect 615 360 655 370
rect 715 640 755 650
rect 715 370 725 640
rect 745 370 755 640
rect 715 360 755 370
rect 795 640 835 650
rect 795 370 805 640
rect 825 370 835 640
rect 795 360 835 370
rect 895 640 935 650
rect 895 370 905 640
rect 925 370 935 640
rect 895 360 935 370
rect 995 640 1035 650
rect 995 370 1005 640
rect 1025 370 1035 640
rect 995 360 1035 370
rect 1075 640 1115 650
rect 1075 370 1085 640
rect 1105 370 1115 640
rect 1075 360 1115 370
rect 1175 640 1215 650
rect 1175 370 1185 640
rect 1205 370 1215 640
rect 1175 360 1215 370
rect 1275 640 1315 650
rect 1275 370 1285 640
rect 1305 370 1315 640
rect 1275 360 1315 370
rect 165 295 185 360
rect 245 295 265 360
rect 445 295 465 360
rect 525 295 545 360
rect 725 295 745 360
rect 805 295 825 360
rect 1005 295 1025 360
rect 1085 295 1105 360
rect -45 285 -5 295
rect -45 15 -35 285
rect -15 15 -5 285
rect -45 5 -5 15
rect 55 285 95 295
rect 55 15 65 285
rect 85 15 95 285
rect 55 5 95 15
rect 155 285 195 295
rect 155 15 165 285
rect 185 15 195 285
rect 155 5 195 15
rect 235 285 275 295
rect 235 15 245 285
rect 265 15 275 285
rect 235 5 275 15
rect 335 285 375 295
rect 335 15 345 285
rect 365 15 375 285
rect 335 5 375 15
rect 435 285 475 295
rect 435 15 445 285
rect 465 15 475 285
rect 435 5 475 15
rect 515 285 555 295
rect 515 15 525 285
rect 545 15 555 285
rect 515 5 555 15
rect 615 285 655 295
rect 615 15 625 285
rect 645 15 655 285
rect 615 5 655 15
rect 715 285 755 295
rect 715 15 725 285
rect 745 15 755 285
rect 715 5 755 15
rect 795 285 835 295
rect 795 15 805 285
rect 825 15 835 285
rect 795 5 835 15
rect 895 285 935 295
rect 895 15 905 285
rect 925 15 935 285
rect 895 5 935 15
rect 995 285 1035 295
rect 995 15 1005 285
rect 1025 15 1035 285
rect 995 5 1035 15
rect 1075 285 1115 295
rect 1075 15 1085 285
rect 1105 15 1115 285
rect 1075 5 1115 15
rect 1175 285 1215 295
rect 1175 15 1185 285
rect 1205 15 1215 285
rect 1175 5 1215 15
rect 1275 285 1315 295
rect 1275 15 1285 285
rect 1305 15 1315 285
rect 1275 5 1315 15
rect 65 -5 85 5
rect 345 -5 365 5
rect 625 -5 645 5
rect 905 -5 925 5
rect 1185 -5 1205 5
rect 5 -25 45 -15
rect 5 -45 15 -25
rect 35 -45 45 -25
rect 5 -55 45 -45
rect 1225 -25 1265 -15
rect 1225 -45 1235 -25
rect 1255 -45 1265 -25
rect 1225 -55 1265 -45
rect 65 -110 85 -90
rect 345 -110 365 -90
rect 625 -110 645 -90
rect 905 -110 925 -90
rect 1185 -110 1205 -90
rect -45 -120 -5 -110
rect -45 -390 -35 -120
rect -15 -390 -5 -120
rect -45 -400 -5 -390
rect 55 -120 95 -110
rect 55 -390 65 -120
rect 85 -390 95 -120
rect 55 -400 95 -390
rect 155 -120 275 -110
rect 155 -390 165 -120
rect 185 -390 245 -120
rect 265 -390 275 -120
rect 155 -400 275 -390
rect 335 -120 375 -110
rect 335 -390 345 -120
rect 365 -390 375 -120
rect 335 -400 375 -390
rect 435 -120 555 -110
rect 435 -390 445 -120
rect 465 -390 525 -120
rect 545 -390 555 -120
rect 435 -400 555 -390
rect 615 -120 655 -110
rect 615 -390 625 -120
rect 645 -390 655 -120
rect 615 -400 655 -390
rect 715 -120 835 -110
rect 715 -390 725 -120
rect 745 -390 805 -120
rect 825 -390 835 -120
rect 715 -400 835 -390
rect 895 -120 935 -110
rect 895 -390 905 -120
rect 925 -390 935 -120
rect 895 -400 935 -390
rect 995 -120 1115 -110
rect 995 -390 1005 -120
rect 1025 -390 1085 -120
rect 1105 -390 1115 -120
rect 995 -400 1115 -390
rect 1175 -120 1215 -110
rect 1175 -390 1185 -120
rect 1205 -390 1215 -120
rect 1175 -400 1215 -390
rect 1275 -120 1315 -110
rect 1275 -390 1285 -120
rect 1305 -390 1315 -120
rect 1275 -400 1315 -390
rect 5 -430 45 -420
rect 5 -450 15 -430
rect 35 -450 45 -430
rect 5 -460 45 -450
rect 1225 -430 1265 -420
rect 1225 -450 1235 -430
rect 1255 -450 1265 -430
rect 1225 -460 1265 -450
<< viali >>
rect -35 1740 -15 2010
rect 165 1740 185 2010
rect 245 1740 265 2010
rect 445 1740 465 2010
rect 525 1740 545 2010
rect 725 1740 745 2010
rect 805 1740 825 2010
rect 1005 1740 1025 2010
rect 1085 1740 1105 2010
rect 1285 1740 1305 2010
rect -35 1270 -15 1540
rect 1285 1270 1305 1540
rect -35 790 -15 1060
rect 165 790 185 1060
rect 245 790 265 1060
rect 445 790 465 1060
rect 525 790 545 1060
rect 725 790 745 1060
rect 805 790 825 1060
rect 1005 790 1025 1060
rect 1085 790 1105 1060
rect 1285 790 1305 1060
rect -35 -390 -15 -120
rect 165 -390 185 -120
rect 245 -390 265 -120
rect 445 -390 465 -120
rect 525 -390 545 -120
rect 725 -390 745 -120
rect 805 -390 825 -120
rect 1005 -390 1025 -120
rect 1085 -390 1105 -120
rect 1285 -390 1305 -120
<< end >>
