magic
tech sky130A
timestamp 1697139793
<< error_p >>
rect -75 782 -55 785
rect -75 518 -72 782
rect -58 518 -55 782
rect -75 515 -55 518
rect 125 782 145 785
rect 125 518 128 782
rect 142 518 145 782
rect 125 515 145 518
rect 305 782 325 785
rect 305 518 308 782
rect 322 518 325 782
rect 305 515 325 518
rect 865 782 885 785
rect 865 518 868 782
rect 882 518 885 782
rect 865 515 885 518
rect 1245 782 1265 785
rect 1245 518 1248 782
rect 1262 518 1265 782
rect 1245 515 1265 518
rect 1425 782 1445 785
rect 1425 518 1428 782
rect 1442 518 1445 782
rect 1425 515 1445 518
<< nmos >>
rect -240 500 -190 800
rect -140 500 -90 800
rect -40 500 10 800
rect 60 500 110 800
rect 160 500 210 800
rect 340 500 390 800
rect 520 500 570 800
rect 620 500 670 800
rect 800 500 850 800
rect 900 500 950 800
rect 1080 500 1130 800
rect 1180 500 1230 800
rect 1360 500 1410 800
rect 1540 500 1590 800
rect 1640 500 1690 800
rect 1740 500 1790 800
rect 1840 500 1890 800
rect 1940 500 1990 800
rect 0 -20 50 280
rect 100 -20 150 280
rect 200 -20 250 280
rect 300 -20 350 280
rect 400 -20 450 280
rect 500 -20 550 280
rect 600 -20 650 280
rect 700 -20 750 280
rect 800 -20 850 280
rect 900 -20 950 280
rect 1000 -20 1050 280
rect 1100 -20 1150 280
rect 1200 -20 1250 280
rect 1300 -20 1350 280
rect 1400 -20 1450 280
rect 1500 -20 1550 280
rect 1600 -20 1650 280
rect 1700 -20 1750 280
<< ndiff >>
rect -290 785 -240 800
rect -290 515 -275 785
rect -255 515 -240 785
rect -290 500 -240 515
rect -190 785 -140 800
rect -190 515 -175 785
rect -155 515 -140 785
rect -190 500 -140 515
rect -90 785 -40 800
rect -90 515 -75 785
rect -55 515 -40 785
rect -90 500 -40 515
rect 10 785 60 800
rect 10 515 25 785
rect 45 515 60 785
rect 10 500 60 515
rect 110 785 160 800
rect 110 515 125 785
rect 145 515 160 785
rect 110 500 160 515
rect 210 785 260 800
rect 210 515 225 785
rect 245 515 260 785
rect 210 500 260 515
rect 290 785 340 800
rect 290 515 305 785
rect 325 515 340 785
rect 290 500 340 515
rect 390 785 440 800
rect 390 515 405 785
rect 425 515 440 785
rect 390 500 440 515
rect 470 785 520 800
rect 470 515 485 785
rect 505 515 520 785
rect 470 500 520 515
rect 570 785 620 800
rect 570 515 585 785
rect 605 515 620 785
rect 570 500 620 515
rect 670 785 720 800
rect 670 515 685 785
rect 705 515 720 785
rect 670 500 720 515
rect 750 785 800 800
rect 750 515 765 785
rect 785 515 800 785
rect 750 500 800 515
rect 850 785 900 800
rect 850 515 865 785
rect 885 515 900 785
rect 850 500 900 515
rect 950 785 1000 800
rect 950 515 965 785
rect 985 515 1000 785
rect 950 500 1000 515
rect 1030 785 1080 800
rect 1030 515 1045 785
rect 1065 515 1080 785
rect 1030 500 1080 515
rect 1130 785 1180 800
rect 1130 515 1145 785
rect 1165 515 1180 785
rect 1130 500 1180 515
rect 1230 785 1280 800
rect 1230 515 1245 785
rect 1265 515 1280 785
rect 1230 500 1280 515
rect 1310 785 1360 800
rect 1310 515 1325 785
rect 1345 515 1360 785
rect 1310 500 1360 515
rect 1410 785 1460 800
rect 1410 515 1425 785
rect 1445 515 1460 785
rect 1410 500 1460 515
rect 1490 785 1540 800
rect 1490 515 1505 785
rect 1525 515 1540 785
rect 1490 500 1540 515
rect 1590 785 1640 800
rect 1590 515 1605 785
rect 1625 515 1640 785
rect 1590 500 1640 515
rect 1690 785 1740 800
rect 1690 515 1705 785
rect 1725 515 1740 785
rect 1690 500 1740 515
rect 1790 785 1840 800
rect 1790 515 1805 785
rect 1825 515 1840 785
rect 1790 500 1840 515
rect 1890 785 1940 800
rect 1890 515 1905 785
rect 1925 515 1940 785
rect 1890 500 1940 515
rect 1990 785 2040 800
rect 1990 515 2005 785
rect 2025 515 2040 785
rect 1990 500 2040 515
rect -50 265 0 280
rect -50 -5 -35 265
rect -15 -5 0 265
rect -50 -20 0 -5
rect 50 265 100 280
rect 50 -5 65 265
rect 85 -5 100 265
rect 50 -20 100 -5
rect 150 265 200 280
rect 150 -5 165 265
rect 185 -5 200 265
rect 150 -20 200 -5
rect 250 265 300 280
rect 250 -5 265 265
rect 285 -5 300 265
rect 250 -20 300 -5
rect 350 265 400 280
rect 350 -5 365 265
rect 385 -5 400 265
rect 350 -20 400 -5
rect 450 265 500 280
rect 450 -5 465 265
rect 485 -5 500 265
rect 450 -20 500 -5
rect 550 265 600 280
rect 550 -5 565 265
rect 585 -5 600 265
rect 550 -20 600 -5
rect 650 265 700 280
rect 650 -5 665 265
rect 685 -5 700 265
rect 650 -20 700 -5
rect 750 265 800 280
rect 750 -5 765 265
rect 785 -5 800 265
rect 750 -20 800 -5
rect 850 265 900 280
rect 850 -5 865 265
rect 885 -5 900 265
rect 850 -20 900 -5
rect 950 265 1000 280
rect 950 -5 965 265
rect 985 -5 1000 265
rect 950 -20 1000 -5
rect 1050 265 1100 280
rect 1050 -5 1065 265
rect 1085 -5 1100 265
rect 1050 -20 1100 -5
rect 1150 265 1200 280
rect 1150 -5 1165 265
rect 1185 -5 1200 265
rect 1150 -20 1200 -5
rect 1250 265 1300 280
rect 1250 -5 1265 265
rect 1285 -5 1300 265
rect 1250 -20 1300 -5
rect 1350 265 1400 280
rect 1350 -5 1365 265
rect 1385 -5 1400 265
rect 1350 -20 1400 -5
rect 1450 265 1500 280
rect 1450 -5 1465 265
rect 1485 -5 1500 265
rect 1450 -20 1500 -5
rect 1550 265 1600 280
rect 1550 -5 1565 265
rect 1585 -5 1600 265
rect 1550 -20 1600 -5
rect 1650 265 1700 280
rect 1650 -5 1665 265
rect 1685 -5 1700 265
rect 1650 -20 1700 -5
rect 1750 265 1800 280
rect 1750 -5 1765 265
rect 1785 -5 1800 265
rect 1750 -20 1800 -5
<< ndiffc >>
rect -275 515 -255 785
rect -175 515 -155 785
rect -75 515 -55 785
rect 25 515 45 785
rect 125 515 145 785
rect 225 515 245 785
rect 305 515 325 785
rect 405 515 425 785
rect 485 515 505 785
rect 585 515 605 785
rect 685 515 705 785
rect 765 515 785 785
rect 865 515 885 785
rect 965 515 985 785
rect 1045 515 1065 785
rect 1145 515 1165 785
rect 1245 515 1265 785
rect 1325 515 1345 785
rect 1425 515 1445 785
rect 1505 515 1525 785
rect 1605 515 1625 785
rect 1705 515 1725 785
rect 1805 515 1825 785
rect 1905 515 1925 785
rect 2005 515 2025 785
rect -35 -5 -15 265
rect 65 -5 85 265
rect 165 -5 185 265
rect 265 -5 285 265
rect 365 -5 385 265
rect 465 -5 485 265
rect 565 -5 585 265
rect 665 -5 685 265
rect 765 -5 785 265
rect 865 -5 885 265
rect 965 -5 985 265
rect 1065 -5 1085 265
rect 1165 -5 1185 265
rect 1265 -5 1285 265
rect 1365 -5 1385 265
rect 1465 -5 1485 265
rect 1565 -5 1585 265
rect 1665 -5 1685 265
rect 1765 -5 1785 265
<< poly >>
rect 695 840 735 850
rect 695 820 705 840
rect 725 820 735 840
rect -240 800 -190 815
rect -140 800 -90 815
rect -40 800 10 815
rect 60 800 110 815
rect 160 800 210 815
rect 340 800 390 815
rect 520 800 570 815
rect 620 800 670 815
rect 695 810 735 820
rect 800 800 850 815
rect 900 800 950 815
rect 1080 800 1130 815
rect 1180 800 1230 815
rect 1360 800 1410 815
rect 1540 800 1590 815
rect 1640 800 1690 815
rect 1740 800 1790 815
rect 1840 800 1890 815
rect 1940 800 1990 815
rect -240 475 -190 500
rect -240 455 -225 475
rect -205 455 -190 475
rect -240 445 -190 455
rect -140 475 -90 500
rect -140 455 -125 475
rect -105 455 -90 475
rect -140 445 -90 455
rect -40 475 10 500
rect -40 455 -25 475
rect -5 455 10 475
rect -40 445 10 455
rect 60 475 110 500
rect 60 455 75 475
rect 95 455 110 475
rect 60 445 110 455
rect 160 475 210 500
rect 160 455 175 475
rect 195 455 210 475
rect 160 445 210 455
rect 340 485 390 500
rect 520 485 570 500
rect 620 485 670 500
rect 800 485 850 500
rect 900 485 950 500
rect 1080 485 1130 500
rect 1180 485 1230 500
rect 1360 485 1410 500
rect 340 475 1410 485
rect 340 455 355 475
rect 375 455 1410 475
rect 340 445 1410 455
rect 1540 475 1590 500
rect 1540 455 1555 475
rect 1575 455 1590 475
rect 1540 445 1590 455
rect 1640 475 1690 500
rect 1640 455 1655 475
rect 1675 455 1690 475
rect 1640 445 1690 455
rect 1740 475 1790 500
rect 1740 455 1755 475
rect 1775 455 1790 475
rect 1740 445 1790 455
rect 1840 475 1890 500
rect 1840 455 1855 475
rect 1875 455 1890 475
rect 1840 445 1890 455
rect 1940 475 1990 500
rect 1940 455 1955 475
rect 1975 455 1990 475
rect 1940 445 1990 455
rect 0 325 50 335
rect 0 305 15 325
rect 35 305 50 325
rect 0 280 50 305
rect 100 325 150 335
rect 100 305 115 325
rect 135 305 150 325
rect 100 280 150 305
rect 200 325 250 335
rect 200 305 215 325
rect 235 305 250 325
rect 200 280 250 305
rect 300 325 350 335
rect 300 305 315 325
rect 335 305 350 325
rect 300 280 350 305
rect 400 325 450 335
rect 400 305 415 325
rect 435 305 450 325
rect 400 280 450 305
rect 500 325 550 335
rect 500 305 515 325
rect 535 305 550 325
rect 500 280 550 305
rect 600 325 650 335
rect 600 305 615 325
rect 635 305 650 325
rect 600 280 650 305
rect 700 325 750 335
rect 700 305 715 325
rect 735 305 750 325
rect 700 280 750 305
rect 800 325 850 335
rect 800 305 815 325
rect 835 305 850 325
rect 800 280 850 305
rect 900 325 950 335
rect 900 305 915 325
rect 935 305 950 325
rect 900 280 950 305
rect 1000 325 1050 335
rect 1000 305 1015 325
rect 1035 305 1050 325
rect 1000 280 1050 305
rect 1100 325 1150 335
rect 1100 305 1115 325
rect 1135 305 1150 325
rect 1100 280 1150 305
rect 1200 325 1250 335
rect 1200 305 1215 325
rect 1235 305 1250 325
rect 1200 280 1250 305
rect 1300 325 1350 335
rect 1300 305 1315 325
rect 1335 305 1350 325
rect 1300 280 1350 305
rect 1400 325 1450 335
rect 1400 305 1415 325
rect 1435 305 1450 325
rect 1400 280 1450 305
rect 1500 325 1550 335
rect 1500 305 1515 325
rect 1535 305 1550 325
rect 1500 280 1550 305
rect 1600 325 1650 335
rect 1600 305 1615 325
rect 1635 305 1650 325
rect 1600 280 1650 305
rect 1700 325 1750 335
rect 1700 305 1715 325
rect 1735 305 1750 325
rect 1700 280 1750 305
rect 0 -35 50 -20
rect 100 -35 150 -20
rect 200 -35 250 -20
rect 300 -35 350 -20
rect 400 -35 450 -20
rect 500 -35 550 -20
rect 600 -35 650 -20
rect 700 -35 750 -20
rect 800 -35 850 -20
rect 900 -35 950 -20
rect 1000 -35 1050 -20
rect 1100 -35 1150 -20
rect 1200 -35 1250 -20
rect 1300 -35 1350 -20
rect 1400 -35 1450 -20
rect 1500 -35 1550 -20
rect 1600 -35 1650 -20
rect 1700 -35 1750 -20
<< polycont >>
rect 705 820 725 840
rect -225 455 -205 475
rect -125 455 -105 475
rect -25 455 -5 475
rect 75 455 95 475
rect 175 455 195 475
rect 355 455 375 475
rect 1555 455 1575 475
rect 1655 455 1675 475
rect 1755 455 1775 475
rect 1855 455 1875 475
rect 1955 455 1975 475
rect 15 305 35 325
rect 115 305 135 325
rect 215 305 235 325
rect 315 305 335 325
rect 415 305 435 325
rect 515 305 535 325
rect 615 305 635 325
rect 715 305 735 325
rect 815 305 835 325
rect 915 305 935 325
rect 1015 305 1035 325
rect 1115 305 1135 325
rect 1215 305 1235 325
rect 1315 305 1335 325
rect 1415 305 1435 325
rect 1515 305 1535 325
rect 1615 305 1635 325
rect 1715 305 1735 325
<< locali >>
rect 415 870 1335 890
rect 415 795 435 870
rect 695 840 735 850
rect 695 820 705 840
rect 725 820 735 840
rect 695 810 735 820
rect 695 795 715 810
rect 765 795 785 870
rect 965 795 985 870
rect 1315 795 1335 870
rect 1490 815 1925 835
rect 1505 795 1525 815
rect 1705 795 1725 815
rect 1905 795 1925 815
rect -285 785 -245 795
rect -285 515 -275 785
rect -255 515 -245 785
rect -285 485 -245 515
rect -185 785 -145 795
rect -185 515 -175 785
rect -155 515 -145 785
rect -185 505 -145 515
rect -85 785 -45 795
rect -85 515 -75 785
rect -55 515 -45 785
rect -85 505 -45 515
rect 15 785 55 795
rect 15 515 25 785
rect 45 515 55 785
rect 15 505 55 515
rect 115 785 155 795
rect 115 515 125 785
rect 145 515 155 785
rect 115 505 155 515
rect 215 785 255 795
rect 215 515 225 785
rect 245 515 255 785
rect 215 505 255 515
rect 295 785 335 795
rect 295 515 305 785
rect 325 515 335 785
rect 295 505 335 515
rect 395 785 435 795
rect 395 515 405 785
rect 425 515 435 785
rect 395 505 435 515
rect 475 785 515 795
rect 475 515 485 785
rect 505 515 515 785
rect 475 505 515 515
rect 575 785 615 795
rect 575 515 585 785
rect 605 515 615 785
rect 575 505 615 515
rect 675 785 715 795
rect 675 515 685 785
rect 705 515 715 785
rect 675 505 715 515
rect 755 785 795 795
rect 755 515 765 785
rect 785 515 795 785
rect 755 505 795 515
rect 855 785 895 795
rect 855 515 865 785
rect 885 515 895 785
rect 855 505 895 515
rect 955 785 995 795
rect 955 515 965 785
rect 985 515 995 785
rect 955 505 995 515
rect 1035 785 1075 795
rect 1035 515 1045 785
rect 1065 515 1075 785
rect 1035 505 1075 515
rect 1135 785 1175 795
rect 1135 515 1145 785
rect 1165 515 1175 785
rect 1135 505 1175 515
rect 1235 785 1275 795
rect 1235 515 1245 785
rect 1265 515 1275 785
rect 1235 505 1275 515
rect 1315 785 1355 795
rect 1315 515 1325 785
rect 1345 515 1355 785
rect 1315 505 1355 515
rect 1415 785 1455 795
rect 1415 515 1425 785
rect 1445 515 1455 785
rect 1415 505 1455 515
rect 1495 785 1535 795
rect 1495 515 1505 785
rect 1525 515 1535 785
rect 1495 505 1535 515
rect 1595 785 1635 795
rect 1595 515 1605 785
rect 1625 515 1635 785
rect 1595 505 1635 515
rect 1695 785 1735 795
rect 1695 515 1705 785
rect 1725 515 1735 785
rect 1695 505 1735 515
rect 1795 785 1835 795
rect 1795 515 1805 785
rect 1825 515 1835 785
rect 1795 505 1835 515
rect 1895 785 1935 795
rect 1895 515 1905 785
rect 1925 515 1935 785
rect 1895 505 1935 515
rect 1995 785 2035 795
rect 1995 515 2005 785
rect 2025 515 2035 785
rect -170 485 -145 505
rect 25 485 45 505
rect 225 485 245 505
rect 495 485 515 505
rect 1035 485 1055 505
rect 1605 485 1625 505
rect 1805 485 1825 505
rect 1995 485 2035 515
rect -285 475 -190 485
rect -285 455 -225 475
rect -205 455 -190 475
rect -285 445 -190 455
rect -170 475 390 485
rect -170 455 -125 475
rect -105 455 -25 475
rect -5 455 75 475
rect 95 455 175 475
rect 195 455 355 475
rect 375 455 390 475
rect 495 465 1055 485
rect 1540 475 1890 485
rect -170 445 390 455
rect 1540 455 1555 475
rect 1575 455 1655 475
rect 1675 455 1755 475
rect 1775 455 1855 475
rect 1875 455 1890 475
rect 1540 445 1890 455
rect 1940 475 2035 485
rect 1940 455 1955 475
rect 1975 455 2035 475
rect 1940 445 2035 455
rect -45 325 50 335
rect -45 305 15 325
rect 35 305 50 325
rect -45 295 50 305
rect 100 325 1650 335
rect 100 305 115 325
rect 135 305 215 325
rect 235 305 315 325
rect 335 305 415 325
rect 435 305 515 325
rect 535 305 615 325
rect 635 305 715 325
rect 735 305 815 325
rect 835 305 915 325
rect 935 305 1015 325
rect 1035 305 1115 325
rect 1135 305 1215 325
rect 1235 305 1315 325
rect 1335 305 1415 325
rect 1435 305 1515 325
rect 1535 305 1615 325
rect 1635 305 1650 325
rect 100 295 1650 305
rect 1700 325 1795 335
rect 1700 305 1715 325
rect 1735 305 1795 325
rect 1700 295 1795 305
rect -45 265 -5 295
rect 165 275 185 295
rect 365 275 385 295
rect 765 275 785 295
rect 965 275 985 295
rect 1365 275 1385 295
rect 1565 275 1585 295
rect -45 -5 -35 265
rect -15 -5 -5 265
rect -45 -15 -5 -5
rect 55 265 95 275
rect 55 -5 65 265
rect 85 -5 95 265
rect 55 -15 95 -5
rect 155 265 195 275
rect 155 -5 165 265
rect 185 -5 195 265
rect 155 -15 195 -5
rect 255 265 295 275
rect 255 -5 265 265
rect 285 -5 295 265
rect 255 -15 295 -5
rect 355 265 395 275
rect 355 -5 365 265
rect 385 -5 395 265
rect 355 -15 395 -5
rect 455 265 495 275
rect 455 -5 465 265
rect 485 -5 495 265
rect 455 -15 495 -5
rect 555 265 595 275
rect 555 -5 565 265
rect 585 -5 595 265
rect 555 -15 595 -5
rect 655 265 695 275
rect 655 -5 665 265
rect 685 -5 695 265
rect 655 -15 695 -5
rect 755 265 795 275
rect 755 -5 765 265
rect 785 -5 795 265
rect 755 -15 795 -5
rect 855 265 895 275
rect 855 -5 865 265
rect 885 -5 895 265
rect 855 -15 895 -5
rect 955 265 995 275
rect 955 -5 965 265
rect 985 -5 995 265
rect 955 -15 995 -5
rect 1055 265 1095 275
rect 1055 -5 1065 265
rect 1085 -5 1095 265
rect 1055 -15 1095 -5
rect 1155 265 1195 275
rect 1155 -5 1165 265
rect 1185 -5 1195 265
rect 1155 -15 1195 -5
rect 1255 265 1295 275
rect 1255 -5 1265 265
rect 1285 -5 1295 265
rect 1255 -15 1295 -5
rect 1355 265 1395 275
rect 1355 -5 1365 265
rect 1385 -5 1395 265
rect 1355 -15 1395 -5
rect 1455 265 1495 275
rect 1455 -5 1465 265
rect 1485 -5 1495 265
rect 1455 -15 1495 -5
rect 1555 265 1595 275
rect 1555 -5 1565 265
rect 1585 -5 1595 265
rect 1555 -15 1595 -5
rect 1655 265 1695 275
rect 1655 -5 1665 265
rect 1685 -5 1695 265
rect 1655 -15 1695 -5
rect 1755 265 1795 295
rect 1755 -5 1765 265
rect 1785 -5 1795 265
rect 1755 -15 1795 -5
rect 65 -35 85 -15
rect 265 -35 285 -15
rect 465 -35 485 -15
rect 665 -35 685 -15
rect 865 -35 885 -15
rect 1065 -35 1085 -15
rect 1265 -35 1285 -15
rect 1465 -35 1485 -15
rect 1665 -35 1685 -15
rect 65 -55 1685 -35
<< viali >>
rect -275 515 -255 785
rect -75 515 -55 785
rect 125 515 145 785
rect 305 515 325 785
rect 865 515 885 785
rect 1245 515 1265 785
rect 1425 515 1445 785
rect 2005 515 2025 785
rect -35 -5 -15 265
rect 565 -5 585 265
rect 1165 -5 1185 265
rect 1765 -5 1785 265
<< metal1 >>
rect -285 785 -245 795
rect 1995 785 2035 795
rect -285 515 -275 785
rect -255 515 -245 785
rect 1995 515 2005 785
rect 2025 515 2035 785
rect -285 505 -245 515
rect 1995 505 2035 515
rect -45 265 -5 275
rect -45 -5 -35 265
rect -15 -5 -5 265
rect -45 -15 -5 -5
rect 555 265 595 275
rect 555 -5 565 265
rect 585 -5 595 265
rect 555 -15 595 -5
rect 1155 265 1195 275
rect 1155 -5 1165 265
rect 1185 -5 1195 265
rect 1155 -15 1195 -5
rect 1755 265 1795 275
rect 1755 -5 1765 265
rect 1785 -5 1795 265
rect 1755 -15 1795 -5
<< labels >>
rlabel locali -170 445 -165 505 5 i
<< end >>
