magic
tech sky130A
timestamp 1694273127
<< nwell >>
rect -120 135 85 375
<< nmos >>
rect 0 0 15 100
<< pmos >>
rect 0 155 15 355
<< ndiff >>
rect -50 85 0 100
rect -50 15 -35 85
rect -15 15 0 85
rect -50 0 0 15
rect 15 85 65 100
rect 15 15 30 85
rect 50 15 65 85
rect 15 0 65 15
<< pdiff >>
rect -50 340 0 355
rect -50 170 -35 340
rect -15 170 0 340
rect -50 155 0 170
rect 15 340 65 355
rect 15 170 30 340
rect 50 170 65 340
rect 15 155 65 170
<< ndiffc >>
rect -35 15 -15 85
rect 30 15 50 85
<< pdiffc >>
rect -35 170 -15 340
rect 30 170 50 340
<< psubdiff >>
rect -100 85 -50 100
rect -100 15 -85 85
rect -65 15 -50 85
rect -100 0 -50 15
<< nsubdiff >>
rect -100 340 -50 355
rect -100 170 -85 340
rect -65 170 -50 340
rect -100 155 -50 170
<< psubdiffcont >>
rect -85 15 -65 85
<< nsubdiffcont >>
rect -85 170 -65 340
<< poly >>
rect 0 355 15 370
rect 0 100 15 155
rect 0 -15 15 0
rect -25 -25 15 -15
rect -25 -45 -15 -25
rect 5 -45 15 -25
rect -25 -55 15 -45
<< polycont >>
rect -15 -45 5 -25
<< locali >>
rect -95 340 -5 350
rect -95 170 -85 340
rect -65 170 -35 340
rect -15 170 -5 340
rect -95 160 -5 170
rect 20 340 60 350
rect 20 170 30 340
rect 50 170 60 340
rect 20 160 60 170
rect 40 95 60 160
rect -95 85 -5 95
rect -95 15 -85 85
rect -65 15 -35 85
rect -15 15 -5 85
rect -95 5 -5 15
rect 20 85 60 95
rect 20 15 30 85
rect 50 15 60 85
rect 20 5 60 15
rect 40 -15 60 5
rect -120 -25 15 -15
rect -120 -35 -15 -25
rect -25 -45 -15 -35
rect 5 -45 15 -25
rect 40 -35 85 -15
rect -25 -55 15 -45
<< viali >>
rect -85 170 -65 340
rect -35 170 -15 340
rect -85 15 -65 85
rect -35 15 -15 85
<< metal1 >>
rect -120 340 85 355
rect -120 170 -85 340
rect -65 170 -35 340
rect -15 170 85 340
rect -120 155 85 170
rect -120 85 85 100
rect -120 15 -85 85
rect -65 15 -35 85
rect -15 15 85 85
rect -120 0 85 15
<< labels >>
rlabel locali -120 -25 -120 -25 7 A
port 1 w
rlabel locali 85 -25 85 -25 3 Y
port 2 e
rlabel metal1 -120 255 -120 255 7 VP
port 3 w
rlabel metal1 -120 50 -120 50 7 VN
port 4 w
<< end >>
