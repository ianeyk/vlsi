magic
tech sky130A
timestamp 1695702519
<< locali >>
rect 2210 660 2230 680
rect 2210 530 2230 550
<< metal1 >>
rect -630 15 -615 30
use flipflop  flipflop_0 ../flipflop
timestamp 1695617576
transform 1 0 -580 0 1 60
box -70 -70 665 900
use flipflop  flipflop_1
timestamp 1695617576
transform 1 0 135 0 1 60
box -70 -70 665 900
use flipflop  flipflop_2
timestamp 1695617576
transform 1 0 850 0 1 60
box -70 -70 665 900
use flipflop  flipflop_3
timestamp 1695617576
transform 1 0 1565 0 1 60
box -70 -70 665 900
<< labels >>
rlabel locali 2230 670 2230 670 3 Q
port 2 e
rlabel locali 2230 540 2230 540 3 Qbar
port 3 e
rlabel metal1 -630 25 -630 25 7 CLK
port 6 w
<< end >>
