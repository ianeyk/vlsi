magic
tech sky130A
timestamp 1695604994
use flipflop_a  flipflop_a_0 ../flipflop
timestamp 1695604286
transform 1 0 105 0 1 80
box -70 -70 665 900
use flipflop_b  flipflop_b_0 ../flipflop
timestamp 1695604286
transform 1 0 820 0 1 80
box -70 -70 665 900
use flipflop_c  flipflop_c_0 ../flipflop
timestamp 1695604286
transform 1 0 1535 0 1 80
box -70 -70 665 900
use flipflop_d  flipflop_d_0 ../flipflop
timestamp 1695604286
transform 1 0 2250 0 1 80
box -70 -70 665 900
<< end >>
