magic
tech sky130A
timestamp 1694264607
<< nwell >>
rect -120 135 200 275
<< nmos >>
rect 10 0 25 100
rect 75 0 90 100
<< pmos >>
rect 0 155 15 255
rect 65 155 80 255
<< ndiff >>
rect -40 85 10 100
rect -40 15 -25 85
rect -5 15 10 85
rect -40 0 10 15
rect 25 0 75 100
rect 90 85 140 100
rect 90 15 105 85
rect 125 15 140 85
rect 90 0 140 15
<< pdiff >>
rect -50 240 0 255
rect -50 170 -35 240
rect -15 170 0 240
rect -50 155 0 170
rect 15 240 65 255
rect 15 170 30 240
rect 50 170 65 240
rect 15 155 65 170
rect 80 240 130 255
rect 80 170 95 240
rect 115 170 130 240
rect 80 155 130 170
<< ndiffc >>
rect -25 15 -5 85
rect 105 15 125 85
<< pdiffc >>
rect -35 170 -15 240
rect 30 170 50 240
rect 95 170 115 240
<< psubdiff >>
rect -120 85 -70 100
rect -120 15 -105 85
rect -85 15 -70 85
rect -120 0 -70 15
rect 140 85 190 100
rect 140 15 155 85
rect 175 15 190 85
rect 140 0 190 15
<< nsubdiff >>
rect -100 240 -50 255
rect -100 170 -85 240
rect -65 170 -50 240
rect -100 155 -50 170
rect 130 240 180 255
rect 130 170 145 240
rect 165 170 180 240
rect 130 155 180 170
<< psubdiffcont >>
rect -105 15 -85 85
rect 155 15 175 85
<< nsubdiffcont >>
rect -85 170 -65 240
rect 145 170 165 240
<< poly >>
rect 0 255 15 270
rect 65 255 80 270
rect 0 130 15 155
rect 65 130 80 155
rect 0 115 25 130
rect 65 115 90 130
rect 10 100 25 115
rect 75 100 90 115
rect 10 -15 25 0
rect -30 -25 25 -15
rect -30 -45 -20 -25
rect 0 -35 25 -25
rect 0 -45 10 -35
rect -30 -55 10 -45
rect 75 -55 90 0
rect 50 -65 90 -55
rect 50 -85 60 -65
rect 80 -85 90 -65
rect 50 -95 90 -85
<< polycont >>
rect -20 -45 0 -25
rect 60 -85 80 -65
<< locali >>
rect -95 240 -5 250
rect -95 170 -85 240
rect -65 170 -35 240
rect -15 170 -5 240
rect -95 160 -5 170
rect 20 240 60 250
rect 20 170 30 240
rect 50 170 60 240
rect 20 160 60 170
rect 85 240 175 250
rect 85 170 95 240
rect 115 170 145 240
rect 165 170 175 240
rect 85 160 175 170
rect 30 95 50 160
rect -115 85 -75 95
rect -115 15 -105 85
rect -85 15 -75 85
rect -115 5 -75 15
rect -35 85 50 95
rect -35 15 -25 85
rect -5 75 50 85
rect -5 15 5 75
rect -35 5 5 15
rect 30 -15 50 75
rect 95 85 185 95
rect 95 15 105 85
rect 125 15 155 85
rect 175 15 185 85
rect 95 5 185 15
rect -120 -25 10 -15
rect -120 -35 -20 -25
rect -30 -45 -20 -35
rect 0 -45 10 -25
rect 30 -35 200 -15
rect -30 -55 10 -45
rect 50 -65 90 -55
rect 50 -75 60 -65
rect -120 -85 60 -75
rect 80 -85 90 -65
rect -120 -95 90 -85
<< viali >>
rect -85 170 -65 240
rect -35 170 -15 240
rect 95 170 115 240
rect 145 170 165 240
rect -105 15 -85 85
rect 105 15 125 85
rect 155 15 175 85
<< metal1 >>
rect -120 240 200 255
rect -120 170 -85 240
rect -65 170 -35 240
rect -15 170 95 240
rect 115 170 145 240
rect 165 170 200 240
rect -120 155 200 170
rect -120 85 200 100
rect -120 15 -105 85
rect -85 15 105 85
rect 125 15 155 85
rect 175 15 200 85
rect -120 0 200 15
<< labels >>
rlabel locali -120 -25 -120 -25 7 A
port 1 w
rlabel locali -120 -85 -120 -85 7 B
port 2 w
rlabel locali 200 -25 200 -25 3 Y
port 3 e
rlabel metal1 -120 205 -120 205 7 VP
port 4 w
rlabel metal1 -120 50 -120 50 7 VN
port 5 w
<< end >>
