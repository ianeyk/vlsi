magic
tech sky130A
timestamp 1695690941
<< locali >>
rect 2210 660 2230 680
rect 2210 530 2230 550
rect -880 490 -860 510
<< metal1 >>
rect -880 530 -865 720
rect -880 300 -865 450
rect -630 15 -615 30
use flipflop  flipflop_0 ../flipflop
timestamp 1695617576
transform 1 0 -580 0 1 60
box -70 -70 665 900
use flipflop  flipflop_1
timestamp 1695617576
transform 1 0 135 0 1 60
box -70 -70 665 900
use flipflop  flipflop_2
timestamp 1695617576
transform 1 0 850 0 1 60
box -70 -70 665 900
use flipflop  flipflop_3
timestamp 1695617576
transform 1 0 1565 0 1 60
box -70 -70 665 900
use inverter  inverter_0
timestamp 1695689994
transform 1 0 -650 0 1 -10
box -230 310 20 755
<< labels >>
rlabel locali 2230 670 2230 670 3 Q
port 2 e
rlabel locali 2230 540 2230 540 3 Qbar
port 3 e
rlabel locali -880 500 -880 500 7 A
port 1 w
rlabel metal1 -880 625 -880 625 7 VP
port 4 w
rlabel metal1 -880 405 -880 405 7 VN
port 5 w
rlabel metal1 -630 25 -630 25 7 CLK
port 6 w
<< end >>
