magic
tech sky130A
timestamp 1695689994
<< nwell >>
rect -230 515 10 755
<< nmos >>
rect -160 365 -145 465
rect -95 365 -80 465
<< pmos >>
rect -160 535 -145 735
rect -95 535 -80 735
<< ndiff >>
rect -210 450 -160 465
rect -210 380 -195 450
rect -175 380 -160 450
rect -210 365 -160 380
rect -145 450 -95 465
rect -145 380 -130 450
rect -110 380 -95 450
rect -145 365 -95 380
rect -80 450 -30 465
rect -80 380 -65 450
rect -45 380 -30 450
rect -80 365 -30 380
<< pdiff >>
rect -210 720 -160 735
rect -210 550 -195 720
rect -175 550 -160 720
rect -210 535 -160 550
rect -145 720 -95 735
rect -145 550 -130 720
rect -110 550 -95 720
rect -145 535 -95 550
rect -80 720 -30 735
rect -80 550 -65 720
rect -45 550 -30 720
rect -80 535 -30 550
<< ndiffc >>
rect -195 380 -175 450
rect -130 380 -110 450
rect -65 380 -45 450
<< pdiffc >>
rect -195 550 -175 720
rect -130 550 -110 720
rect -65 550 -45 720
<< poly >>
rect -160 735 -145 750
rect -95 735 -80 750
rect -160 520 -145 535
rect -185 510 -145 520
rect -185 490 -175 510
rect -155 490 -145 510
rect -185 480 -145 490
rect -160 465 -145 480
rect -95 465 -80 535
rect -160 350 -145 365
rect -95 350 -80 365
rect -120 340 -80 350
rect -120 320 -110 340
rect -90 320 -80 340
rect -120 310 -80 320
<< polycont >>
rect -175 490 -155 510
rect -110 320 -90 340
<< locali >>
rect -205 720 -165 730
rect -205 550 -195 720
rect -175 550 -165 720
rect -205 540 -165 550
rect -140 720 -100 730
rect -140 550 -130 720
rect -110 550 -100 720
rect -140 540 -100 550
rect -75 720 -35 730
rect -75 550 -65 720
rect -45 690 -35 720
rect -45 670 20 690
rect -45 550 -35 670
rect -75 540 -35 550
rect -230 510 -145 520
rect -230 500 -175 510
rect -185 490 -175 500
rect -155 490 -145 510
rect -185 480 -145 490
rect -55 460 -35 540
rect -205 450 -165 460
rect -205 380 -195 450
rect -175 380 -165 450
rect -205 370 -165 380
rect -140 450 -100 460
rect -140 380 -130 450
rect -110 380 -100 450
rect -140 370 -100 380
rect -75 450 -35 460
rect -75 380 -65 450
rect -45 380 -35 450
rect -75 370 -35 380
rect -15 540 20 560
rect -185 350 -165 370
rect -15 350 5 540
rect -185 340 5 350
rect -185 330 -110 340
rect -120 320 -110 330
rect -90 330 5 340
rect -90 320 -80 330
rect -120 310 -80 320
<< viali >>
rect -130 550 -110 720
rect -130 380 -110 450
<< metal1 >>
rect -230 720 20 730
rect -230 550 -130 720
rect -110 550 20 720
rect -230 540 20 550
rect -230 450 20 460
rect -230 380 -130 450
rect -110 380 20 450
rect -230 310 20 380
<< end >>
