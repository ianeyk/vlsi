magic
tech sky130A
timestamp 1697029401
<< error_p >>
rect -35 2047 -15 2050
rect -35 1783 -32 2047
rect -18 1783 -15 2047
rect -35 1780 -15 1783
rect 165 2047 185 2050
rect 165 1783 168 2047
rect 182 1783 185 2047
rect 165 1780 185 1783
rect 245 2047 265 2050
rect 245 1783 248 2047
rect 262 1783 265 2047
rect 245 1780 265 1783
rect 445 2047 465 2050
rect 445 1783 448 2047
rect 462 1783 465 2047
rect 445 1780 465 1783
rect 525 2047 545 2050
rect 525 1783 528 2047
rect 542 1783 545 2047
rect 525 1780 545 1783
rect 725 2047 745 2050
rect 725 1783 728 2047
rect 742 1783 745 2047
rect 725 1780 745 1783
rect 805 2047 825 2050
rect 805 1783 808 2047
rect 822 1783 825 2047
rect 805 1780 825 1783
rect 1005 2047 1025 2050
rect 1005 1783 1008 2047
rect 1022 1783 1025 2047
rect 1005 1780 1025 1783
rect 1085 2047 1105 2050
rect 1085 1783 1088 2047
rect 1102 1783 1105 2047
rect 1085 1780 1105 1783
rect 1285 2047 1305 2050
rect 1285 1783 1288 2047
rect 1302 1783 1305 2047
rect 1285 1780 1305 1783
rect -35 1577 -15 1580
rect -35 1313 -32 1577
rect -18 1313 -15 1577
rect -35 1310 -15 1313
rect 1285 1577 1305 1580
rect 1285 1313 1288 1577
rect 1302 1313 1305 1577
rect 1285 1310 1305 1313
rect -35 1097 -15 1100
rect -35 833 -32 1097
rect -18 833 -15 1097
rect -35 830 -15 833
rect 165 1097 185 1100
rect 165 833 168 1097
rect 182 833 185 1097
rect 165 830 185 833
rect 245 1097 265 1100
rect 245 833 248 1097
rect 262 833 265 1097
rect 245 830 265 833
rect 445 1097 465 1100
rect 445 833 448 1097
rect 462 833 465 1097
rect 445 830 465 833
rect 525 1097 545 1100
rect 525 833 528 1097
rect 542 833 545 1097
rect 525 830 545 833
rect 725 1097 745 1100
rect 725 833 728 1097
rect 742 833 745 1097
rect 725 830 745 833
rect 805 1097 825 1100
rect 805 833 808 1097
rect 822 833 825 1097
rect 805 830 825 833
rect 1005 1097 1025 1100
rect 1005 833 1008 1097
rect 1022 833 1025 1097
rect 1005 830 1025 833
rect 1085 1097 1105 1100
rect 1085 833 1088 1097
rect 1102 833 1105 1097
rect 1085 830 1105 833
rect 1285 1097 1305 1100
rect 1285 833 1288 1097
rect 1302 833 1305 1097
rect 1285 830 1305 833
rect -35 -123 -15 -120
rect -35 -387 -32 -123
rect -18 -387 -15 -123
rect -35 -390 -15 -387
rect 165 -123 185 -120
rect 165 -387 168 -123
rect 182 -387 185 -123
rect 165 -390 185 -387
rect 245 -123 265 -120
rect 245 -387 248 -123
rect 262 -387 265 -123
rect 245 -390 265 -387
rect 445 -123 465 -120
rect 445 -387 448 -123
rect 462 -387 465 -123
rect 445 -390 465 -387
rect 525 -123 545 -120
rect 525 -387 528 -123
rect 542 -387 545 -123
rect 525 -390 545 -387
rect 725 -123 745 -120
rect 725 -387 728 -123
rect 742 -387 745 -123
rect 725 -390 745 -387
rect 805 -123 825 -120
rect 805 -387 808 -123
rect 822 -387 825 -123
rect 805 -390 825 -387
rect 1005 -123 1025 -120
rect 1005 -387 1008 -123
rect 1022 -387 1025 -123
rect 1005 -390 1025 -387
rect 1085 -123 1105 -120
rect 1085 -387 1088 -123
rect 1102 -387 1105 -123
rect 1085 -390 1105 -387
rect 1285 -123 1305 -120
rect 1285 -387 1288 -123
rect 1302 -387 1305 -123
rect 1285 -390 1305 -387
<< nwell >>
rect -70 375 1340 1135
<< nmos >>
rect 0 1765 50 2065
rect 100 1765 150 2065
rect 280 1765 330 2065
rect 380 1765 430 2065
rect 560 1765 610 2065
rect 660 1765 710 2065
rect 840 1765 890 2065
rect 940 1765 990 2065
rect 1120 1765 1170 2065
rect 1220 1765 1270 2065
rect 0 1295 50 1595
rect 100 1295 150 1595
rect 280 1295 330 1595
rect 380 1295 430 1595
rect 560 1295 610 1595
rect 660 1295 710 1595
rect 840 1295 890 1595
rect 940 1295 990 1595
rect 1120 1295 1170 1595
rect 1220 1295 1270 1595
rect 0 0 50 300
rect 100 0 150 300
rect 280 0 330 300
rect 380 0 430 300
rect 560 0 610 300
rect 660 0 710 300
rect 840 0 890 300
rect 940 0 990 300
rect 1120 0 1170 300
rect 1220 0 1270 300
rect 0 -405 50 -105
rect 100 -405 150 -105
rect 280 -405 330 -105
rect 380 -405 430 -105
rect 560 -405 610 -105
rect 660 -405 710 -105
rect 840 -405 890 -105
rect 940 -405 990 -105
rect 1120 -405 1170 -105
rect 1220 -405 1270 -105
<< pmos >>
rect 0 815 50 1115
rect 100 815 150 1115
rect 280 815 330 1115
rect 380 815 430 1115
rect 560 815 610 1115
rect 660 815 710 1115
rect 840 815 890 1115
rect 940 815 990 1115
rect 1120 815 1170 1115
rect 1220 815 1270 1115
rect 0 395 50 695
rect 100 395 150 695
rect 280 395 330 695
rect 380 395 430 695
rect 560 395 610 695
rect 660 395 710 695
rect 840 395 890 695
rect 940 395 990 695
rect 1120 395 1170 695
rect 1220 395 1270 695
<< ndiff >>
rect -50 2050 0 2065
rect -50 1780 -35 2050
rect -15 1780 0 2050
rect -50 1765 0 1780
rect 50 2050 100 2065
rect 50 1780 65 2050
rect 85 1780 100 2050
rect 50 1765 100 1780
rect 150 2050 200 2065
rect 150 1780 165 2050
rect 185 1780 200 2050
rect 150 1765 200 1780
rect 230 2050 280 2065
rect 230 1780 245 2050
rect 265 1780 280 2050
rect 230 1765 280 1780
rect 330 2050 380 2065
rect 330 1780 345 2050
rect 365 1780 380 2050
rect 330 1765 380 1780
rect 430 2050 480 2065
rect 430 1780 445 2050
rect 465 1780 480 2050
rect 430 1765 480 1780
rect 510 2050 560 2065
rect 510 1780 525 2050
rect 545 1780 560 2050
rect 510 1765 560 1780
rect 610 2050 660 2065
rect 610 1780 625 2050
rect 645 1780 660 2050
rect 610 1765 660 1780
rect 710 2050 760 2065
rect 710 1780 725 2050
rect 745 1780 760 2050
rect 710 1765 760 1780
rect 790 2050 840 2065
rect 790 1780 805 2050
rect 825 1780 840 2050
rect 790 1765 840 1780
rect 890 2050 940 2065
rect 890 1780 905 2050
rect 925 1780 940 2050
rect 890 1765 940 1780
rect 990 2050 1040 2065
rect 990 1780 1005 2050
rect 1025 1780 1040 2050
rect 990 1765 1040 1780
rect 1070 2050 1120 2065
rect 1070 1780 1085 2050
rect 1105 1780 1120 2050
rect 1070 1765 1120 1780
rect 1170 2050 1220 2065
rect 1170 1780 1185 2050
rect 1205 1780 1220 2050
rect 1170 1765 1220 1780
rect 1270 2050 1320 2065
rect 1270 1780 1285 2050
rect 1305 1780 1320 2050
rect 1270 1765 1320 1780
rect -50 1580 0 1595
rect -50 1310 -35 1580
rect -15 1310 0 1580
rect -50 1295 0 1310
rect 50 1580 100 1595
rect 50 1310 65 1580
rect 85 1310 100 1580
rect 50 1295 100 1310
rect 150 1580 200 1595
rect 150 1310 165 1580
rect 185 1310 200 1580
rect 150 1295 200 1310
rect 230 1580 280 1595
rect 230 1310 245 1580
rect 265 1310 280 1580
rect 230 1295 280 1310
rect 330 1580 380 1595
rect 330 1310 345 1580
rect 365 1310 380 1580
rect 330 1295 380 1310
rect 430 1580 480 1595
rect 430 1310 445 1580
rect 465 1310 480 1580
rect 430 1295 480 1310
rect 510 1580 560 1595
rect 510 1310 525 1580
rect 545 1310 560 1580
rect 510 1295 560 1310
rect 610 1580 660 1595
rect 610 1310 625 1580
rect 645 1310 660 1580
rect 610 1295 660 1310
rect 710 1580 760 1595
rect 710 1310 725 1580
rect 745 1310 760 1580
rect 710 1295 760 1310
rect 790 1580 840 1595
rect 790 1310 805 1580
rect 825 1310 840 1580
rect 790 1295 840 1310
rect 890 1580 940 1595
rect 890 1310 905 1580
rect 925 1310 940 1580
rect 890 1295 940 1310
rect 990 1580 1040 1595
rect 990 1310 1005 1580
rect 1025 1310 1040 1580
rect 990 1295 1040 1310
rect 1070 1580 1120 1595
rect 1070 1310 1085 1580
rect 1105 1310 1120 1580
rect 1070 1295 1120 1310
rect 1170 1580 1220 1595
rect 1170 1310 1185 1580
rect 1205 1310 1220 1580
rect 1170 1295 1220 1310
rect 1270 1580 1320 1595
rect 1270 1310 1285 1580
rect 1305 1310 1320 1580
rect 1270 1295 1320 1310
rect -50 285 0 300
rect -50 15 -35 285
rect -15 15 0 285
rect -50 0 0 15
rect 50 285 100 300
rect 50 15 65 285
rect 85 15 100 285
rect 50 0 100 15
rect 150 285 200 300
rect 150 15 165 285
rect 185 15 200 285
rect 150 0 200 15
rect 230 285 280 300
rect 230 15 245 285
rect 265 15 280 285
rect 230 0 280 15
rect 330 285 380 300
rect 330 15 345 285
rect 365 15 380 285
rect 330 0 380 15
rect 430 285 480 300
rect 430 15 445 285
rect 465 15 480 285
rect 430 0 480 15
rect 510 285 560 300
rect 510 15 525 285
rect 545 15 560 285
rect 510 0 560 15
rect 610 285 660 300
rect 610 15 625 285
rect 645 15 660 285
rect 610 0 660 15
rect 710 285 760 300
rect 710 15 725 285
rect 745 15 760 285
rect 710 0 760 15
rect 790 285 840 300
rect 790 15 805 285
rect 825 15 840 285
rect 790 0 840 15
rect 890 285 940 300
rect 890 15 905 285
rect 925 15 940 285
rect 890 0 940 15
rect 990 285 1040 300
rect 990 15 1005 285
rect 1025 15 1040 285
rect 990 0 1040 15
rect 1070 285 1120 300
rect 1070 15 1085 285
rect 1105 15 1120 285
rect 1070 0 1120 15
rect 1170 285 1220 300
rect 1170 15 1185 285
rect 1205 15 1220 285
rect 1170 0 1220 15
rect 1270 285 1320 300
rect 1270 15 1285 285
rect 1305 15 1320 285
rect 1270 0 1320 15
rect -50 -120 0 -105
rect -50 -390 -35 -120
rect -15 -390 0 -120
rect -50 -405 0 -390
rect 50 -120 100 -105
rect 50 -390 65 -120
rect 85 -390 100 -120
rect 50 -405 100 -390
rect 150 -120 200 -105
rect 150 -390 165 -120
rect 185 -390 200 -120
rect 150 -405 200 -390
rect 230 -120 280 -105
rect 230 -390 245 -120
rect 265 -390 280 -120
rect 230 -405 280 -390
rect 330 -120 380 -105
rect 330 -390 345 -120
rect 365 -390 380 -120
rect 330 -405 380 -390
rect 430 -120 480 -105
rect 430 -390 445 -120
rect 465 -390 480 -120
rect 430 -405 480 -390
rect 510 -120 560 -105
rect 510 -390 525 -120
rect 545 -390 560 -120
rect 510 -405 560 -390
rect 610 -120 660 -105
rect 610 -390 625 -120
rect 645 -390 660 -120
rect 610 -405 660 -390
rect 710 -120 760 -105
rect 710 -390 725 -120
rect 745 -390 760 -120
rect 710 -405 760 -390
rect 790 -120 840 -105
rect 790 -390 805 -120
rect 825 -390 840 -120
rect 790 -405 840 -390
rect 890 -120 940 -105
rect 890 -390 905 -120
rect 925 -390 940 -120
rect 890 -405 940 -390
rect 990 -120 1040 -105
rect 990 -390 1005 -120
rect 1025 -390 1040 -120
rect 990 -405 1040 -390
rect 1070 -120 1120 -105
rect 1070 -390 1085 -120
rect 1105 -390 1120 -120
rect 1070 -405 1120 -390
rect 1170 -120 1220 -105
rect 1170 -390 1185 -120
rect 1205 -390 1220 -120
rect 1170 -405 1220 -390
rect 1270 -120 1320 -105
rect 1270 -390 1285 -120
rect 1305 -390 1320 -120
rect 1270 -405 1320 -390
<< pdiff >>
rect -50 1100 0 1115
rect -50 830 -35 1100
rect -15 830 0 1100
rect -50 815 0 830
rect 50 1100 100 1115
rect 50 830 65 1100
rect 85 830 100 1100
rect 50 815 100 830
rect 150 1100 200 1115
rect 150 830 165 1100
rect 185 830 200 1100
rect 150 815 200 830
rect 230 1100 280 1115
rect 230 830 245 1100
rect 265 830 280 1100
rect 230 815 280 830
rect 330 1100 380 1115
rect 330 830 345 1100
rect 365 830 380 1100
rect 330 815 380 830
rect 430 1100 480 1115
rect 430 830 445 1100
rect 465 830 480 1100
rect 430 815 480 830
rect 510 1100 560 1115
rect 510 830 525 1100
rect 545 830 560 1100
rect 510 815 560 830
rect 610 1100 660 1115
rect 610 830 625 1100
rect 645 830 660 1100
rect 610 815 660 830
rect 710 1100 760 1115
rect 710 830 725 1100
rect 745 830 760 1100
rect 710 815 760 830
rect 790 1100 840 1115
rect 790 830 805 1100
rect 825 830 840 1100
rect 790 815 840 830
rect 890 1100 940 1115
rect 890 830 905 1100
rect 925 830 940 1100
rect 890 815 940 830
rect 990 1100 1040 1115
rect 990 830 1005 1100
rect 1025 830 1040 1100
rect 990 815 1040 830
rect 1070 1100 1120 1115
rect 1070 830 1085 1100
rect 1105 830 1120 1100
rect 1070 815 1120 830
rect 1170 1100 1220 1115
rect 1170 830 1185 1100
rect 1205 830 1220 1100
rect 1170 815 1220 830
rect 1270 1100 1320 1115
rect 1270 830 1285 1100
rect 1305 830 1320 1100
rect 1270 815 1320 830
rect -50 680 0 695
rect -50 410 -35 680
rect -15 410 0 680
rect -50 395 0 410
rect 50 680 100 695
rect 50 410 65 680
rect 85 410 100 680
rect 50 395 100 410
rect 150 680 200 695
rect 150 410 165 680
rect 185 410 200 680
rect 150 395 200 410
rect 230 680 280 695
rect 230 410 245 680
rect 265 410 280 680
rect 230 395 280 410
rect 330 680 380 695
rect 330 410 345 680
rect 365 410 380 680
rect 330 395 380 410
rect 430 680 480 695
rect 430 410 445 680
rect 465 410 480 680
rect 430 395 480 410
rect 510 680 560 695
rect 510 410 525 680
rect 545 410 560 680
rect 510 395 560 410
rect 610 680 660 695
rect 610 410 625 680
rect 645 410 660 680
rect 610 395 660 410
rect 710 680 760 695
rect 710 410 725 680
rect 745 410 760 680
rect 710 395 760 410
rect 790 680 840 695
rect 790 410 805 680
rect 825 410 840 680
rect 790 395 840 410
rect 890 680 940 695
rect 890 410 905 680
rect 925 410 940 680
rect 890 395 940 410
rect 990 680 1040 695
rect 990 410 1005 680
rect 1025 410 1040 680
rect 990 395 1040 410
rect 1070 680 1120 695
rect 1070 410 1085 680
rect 1105 410 1120 680
rect 1070 395 1120 410
rect 1170 680 1220 695
rect 1170 410 1185 680
rect 1205 410 1220 680
rect 1170 395 1220 410
rect 1270 680 1320 695
rect 1270 410 1285 680
rect 1305 410 1320 680
rect 1270 395 1320 410
<< ndiffc >>
rect -35 1780 -15 2050
rect 65 1780 85 2050
rect 165 1780 185 2050
rect 245 1780 265 2050
rect 345 1780 365 2050
rect 445 1780 465 2050
rect 525 1780 545 2050
rect 625 1780 645 2050
rect 725 1780 745 2050
rect 805 1780 825 2050
rect 905 1780 925 2050
rect 1005 1780 1025 2050
rect 1085 1780 1105 2050
rect 1185 1780 1205 2050
rect 1285 1780 1305 2050
rect -35 1310 -15 1580
rect 65 1310 85 1580
rect 165 1310 185 1580
rect 245 1310 265 1580
rect 345 1310 365 1580
rect 445 1310 465 1580
rect 525 1310 545 1580
rect 625 1310 645 1580
rect 725 1310 745 1580
rect 805 1310 825 1580
rect 905 1310 925 1580
rect 1005 1310 1025 1580
rect 1085 1310 1105 1580
rect 1185 1310 1205 1580
rect 1285 1310 1305 1580
rect -35 15 -15 285
rect 65 15 85 285
rect 165 15 185 285
rect 245 15 265 285
rect 345 15 365 285
rect 445 15 465 285
rect 525 15 545 285
rect 625 15 645 285
rect 725 15 745 285
rect 805 15 825 285
rect 905 15 925 285
rect 1005 15 1025 285
rect 1085 15 1105 285
rect 1185 15 1205 285
rect 1285 15 1305 285
rect -35 -390 -15 -120
rect 65 -390 85 -120
rect 165 -390 185 -120
rect 245 -390 265 -120
rect 345 -390 365 -120
rect 445 -390 465 -120
rect 525 -390 545 -120
rect 625 -390 645 -120
rect 725 -390 745 -120
rect 805 -390 825 -120
rect 905 -390 925 -120
rect 1005 -390 1025 -120
rect 1085 -390 1105 -120
rect 1185 -390 1205 -120
rect 1285 -390 1305 -120
<< pdiffc >>
rect -35 830 -15 1100
rect 65 830 85 1100
rect 165 830 185 1100
rect 245 830 265 1100
rect 345 830 365 1100
rect 445 830 465 1100
rect 525 830 545 1100
rect 625 830 645 1100
rect 725 830 745 1100
rect 805 830 825 1100
rect 905 830 925 1100
rect 1005 830 1025 1100
rect 1085 830 1105 1100
rect 1185 830 1205 1100
rect 1285 830 1305 1100
rect -35 410 -15 680
rect 65 410 85 680
rect 165 410 185 680
rect 245 410 265 680
rect 345 410 365 680
rect 445 410 465 680
rect 525 410 545 680
rect 625 410 645 680
rect 725 410 745 680
rect 805 410 825 680
rect 905 410 925 680
rect 1005 410 1025 680
rect 1085 410 1105 680
rect 1185 410 1205 680
rect 1285 410 1305 680
<< poly >>
rect 0 2110 50 2120
rect 0 2090 15 2110
rect 35 2090 50 2110
rect 0 2065 50 2090
rect 100 2080 1170 2130
rect 100 2065 150 2080
rect 280 2065 330 2080
rect 380 2065 430 2080
rect 560 2065 610 2080
rect 660 2065 710 2080
rect 840 2065 890 2080
rect 940 2065 990 2080
rect 1120 2065 1170 2080
rect 1220 2110 1270 2120
rect 1220 2090 1235 2110
rect 1255 2090 1270 2110
rect 1220 2065 1270 2090
rect 0 1750 50 1765
rect 100 1750 150 1765
rect 280 1750 330 1765
rect 380 1750 430 1765
rect 560 1750 610 1765
rect 660 1750 710 1765
rect 840 1750 890 1765
rect 940 1750 990 1765
rect 1120 1750 1170 1765
rect 1220 1750 1270 1765
rect -50 1685 125 1725
rect -50 1675 990 1685
rect 0 1640 50 1650
rect 0 1620 15 1640
rect 35 1620 50 1640
rect 75 1635 990 1675
rect 0 1595 50 1620
rect 100 1595 150 1610
rect 280 1595 330 1635
rect 380 1595 430 1635
rect 560 1595 610 1610
rect 660 1595 710 1610
rect 840 1595 890 1635
rect 940 1595 990 1635
rect 1220 1640 1270 1650
rect 1220 1620 1235 1640
rect 1255 1620 1270 1640
rect 1120 1595 1170 1610
rect 1220 1595 1270 1620
rect 0 1280 50 1295
rect 100 1255 150 1295
rect 280 1280 330 1295
rect 380 1280 430 1295
rect 560 1255 610 1295
rect 660 1255 710 1295
rect 840 1280 890 1295
rect 940 1280 990 1295
rect 1120 1255 1170 1295
rect 1220 1280 1270 1295
rect -50 1205 1170 1255
rect 0 1160 50 1170
rect 0 1140 15 1160
rect 35 1140 50 1160
rect 0 1115 50 1140
rect 100 1130 1170 1180
rect 100 1115 150 1130
rect 280 1115 330 1130
rect 380 1115 430 1130
rect 560 1115 610 1130
rect 660 1115 710 1130
rect 840 1115 890 1130
rect 940 1115 990 1130
rect 1120 1115 1170 1130
rect 1220 1160 1270 1170
rect 1220 1140 1235 1160
rect 1255 1140 1270 1160
rect 1220 1115 1270 1140
rect 0 800 50 815
rect 100 800 150 815
rect 280 800 330 815
rect 380 800 430 815
rect 560 800 610 815
rect 660 800 710 815
rect 840 800 890 815
rect 940 800 990 815
rect 1120 800 1170 815
rect 1220 800 1270 815
rect 0 740 50 750
rect 0 720 15 740
rect 35 720 50 740
rect 0 695 50 720
rect 100 710 1170 760
rect 100 695 150 710
rect 280 695 330 710
rect 380 695 430 710
rect 560 695 610 710
rect 660 695 710 710
rect 840 695 890 710
rect 940 695 990 710
rect 1120 695 1170 710
rect 1220 740 1270 750
rect 1220 720 1235 740
rect 1255 720 1270 740
rect 1220 695 1270 720
rect 0 380 50 395
rect 100 380 150 395
rect 280 380 330 395
rect 380 380 430 395
rect 560 380 610 395
rect 660 380 710 395
rect 840 380 890 395
rect 940 380 990 395
rect 1120 380 1170 395
rect 1220 380 1270 395
rect 475 345 805 355
rect 475 325 485 345
rect 505 340 775 345
rect 505 325 515 340
rect 475 315 515 325
rect 765 325 775 340
rect 795 325 805 345
rect 765 315 805 325
rect 0 300 50 315
rect 100 300 150 315
rect 280 300 330 315
rect 380 300 430 315
rect 560 300 610 315
rect 660 300 710 315
rect 840 300 890 315
rect 940 300 990 315
rect 1120 300 1170 315
rect 1220 300 1270 315
rect 0 -25 50 0
rect 0 -45 15 -25
rect 35 -45 50 -25
rect 0 -55 50 -45
rect 100 -15 150 0
rect 280 -15 330 0
rect 380 -15 430 0
rect 560 -15 610 0
rect 660 -15 710 0
rect 840 -15 890 0
rect 940 -15 990 0
rect 1120 -15 1170 0
rect 100 -65 1170 -15
rect 1220 -25 1270 0
rect 1220 -45 1235 -25
rect 1255 -45 1270 -25
rect 1220 -55 1270 -45
rect 0 -105 50 -90
rect 100 -105 150 -90
rect 280 -105 330 -90
rect 380 -105 430 -90
rect 560 -105 610 -90
rect 660 -105 710 -90
rect 840 -105 890 -90
rect 940 -105 990 -90
rect 1120 -105 1170 -90
rect 1220 -105 1270 -90
rect 0 -430 50 -405
rect 0 -450 15 -430
rect 35 -450 50 -430
rect 0 -460 50 -450
rect 100 -420 150 -405
rect 280 -420 330 -405
rect 380 -420 430 -405
rect 560 -420 610 -405
rect 660 -420 710 -405
rect 840 -420 890 -405
rect 940 -420 990 -405
rect 1120 -420 1170 -405
rect 100 -470 1170 -420
rect 1220 -430 1270 -405
rect 1220 -450 1235 -430
rect 1255 -450 1270 -430
rect 1220 -460 1270 -450
<< polycont >>
rect 15 2090 35 2110
rect 1235 2090 1255 2110
rect 15 1620 35 1640
rect 1235 1620 1255 1640
rect 15 1140 35 1160
rect 1235 1140 1255 1160
rect 15 720 35 740
rect 1235 720 1255 740
rect 485 325 505 345
rect 775 325 795 345
rect 15 -45 35 -25
rect 1235 -45 1255 -25
rect 15 -450 35 -430
rect 1235 -450 1255 -430
<< locali >>
rect 5 2110 45 2120
rect 5 2090 15 2110
rect 35 2090 45 2110
rect 5 2080 45 2090
rect 1225 2110 1265 2120
rect 1225 2090 1235 2110
rect 1255 2090 1265 2110
rect 1225 2080 1265 2090
rect -45 2050 -5 2060
rect -45 1780 -35 2050
rect -15 1780 -5 2050
rect -45 1770 -5 1780
rect 55 2050 95 2060
rect 55 1780 65 2050
rect 85 1780 95 2050
rect 55 1770 95 1780
rect 155 2050 275 2060
rect 155 1780 165 2050
rect 185 1780 245 2050
rect 265 1780 275 2050
rect 155 1770 275 1780
rect 335 2050 375 2060
rect 335 1780 345 2050
rect 365 1780 375 2050
rect 335 1770 375 1780
rect 435 2050 555 2060
rect 435 1780 445 2050
rect 465 1780 525 2050
rect 545 1780 555 2050
rect 435 1770 555 1780
rect 615 2050 655 2060
rect 615 1780 625 2050
rect 645 1780 655 2050
rect 615 1770 655 1780
rect 715 2050 835 2060
rect 715 1780 725 2050
rect 745 1780 805 2050
rect 825 1780 835 2050
rect 715 1770 835 1780
rect 895 2050 935 2060
rect 895 1780 905 2050
rect 925 1780 935 2050
rect 895 1770 935 1780
rect 995 2050 1115 2060
rect 995 1780 1005 2050
rect 1025 1780 1085 2050
rect 1105 1780 1115 2050
rect 995 1770 1115 1780
rect 1175 2050 1215 2060
rect 1175 1780 1185 2050
rect 1205 1780 1215 2050
rect 1175 1770 1215 1780
rect 1275 2050 1315 2060
rect 1275 1780 1285 2050
rect 1305 1780 1315 2050
rect 1275 1770 1315 1780
rect 75 1690 95 1770
rect 345 1690 365 1770
rect 625 1690 645 1770
rect 905 1690 925 1770
rect 1175 1690 1195 1770
rect 75 1670 1195 1690
rect 5 1640 45 1650
rect 5 1620 15 1640
rect 35 1620 45 1640
rect 5 1610 45 1620
rect 205 1590 225 1670
rect 485 1590 505 1670
rect 765 1590 785 1670
rect 1045 1590 1065 1670
rect 1225 1640 1265 1650
rect 1225 1620 1235 1640
rect 1255 1620 1265 1640
rect 1225 1610 1265 1620
rect -45 1580 -5 1590
rect -45 1310 -35 1580
rect -15 1310 -5 1580
rect -45 1300 -5 1310
rect 55 1580 95 1590
rect 55 1310 65 1580
rect 85 1310 95 1580
rect 55 1300 95 1310
rect 155 1580 275 1590
rect 155 1310 165 1580
rect 185 1310 245 1580
rect 265 1310 275 1580
rect 155 1300 275 1310
rect 335 1580 375 1590
rect 335 1310 345 1580
rect 365 1310 375 1580
rect 335 1300 375 1310
rect 435 1580 555 1590
rect 435 1310 445 1580
rect 465 1310 525 1580
rect 545 1310 555 1580
rect 435 1300 555 1310
rect 615 1580 655 1590
rect 615 1310 625 1580
rect 645 1310 655 1580
rect 615 1300 655 1310
rect 715 1580 835 1590
rect 715 1310 725 1580
rect 745 1310 805 1580
rect 825 1310 835 1580
rect 715 1300 835 1310
rect 895 1580 935 1590
rect 895 1310 905 1580
rect 925 1310 935 1580
rect 895 1300 935 1310
rect 995 1580 1115 1590
rect 995 1310 1005 1580
rect 1025 1310 1085 1580
rect 1105 1310 1115 1580
rect 995 1300 1115 1310
rect 1175 1580 1215 1590
rect 1175 1310 1185 1580
rect 1205 1310 1215 1580
rect 1175 1300 1215 1310
rect 1275 1580 1315 1590
rect 1275 1310 1285 1580
rect 1305 1310 1315 1580
rect 1275 1300 1315 1310
rect 5 1160 45 1170
rect 5 1140 15 1160
rect 35 1140 45 1160
rect 5 1130 45 1140
rect 65 1110 85 1300
rect 345 1110 365 1300
rect 625 1110 645 1300
rect 905 1110 925 1300
rect 1185 1110 1205 1300
rect 1225 1160 1265 1170
rect 1225 1140 1235 1160
rect 1255 1140 1265 1160
rect 1225 1130 1265 1140
rect -45 1100 -5 1110
rect -45 830 -35 1100
rect -15 830 -5 1100
rect -45 820 -5 830
rect 55 1100 95 1110
rect 55 830 65 1100
rect 85 830 95 1100
rect 55 820 95 830
rect 155 1100 275 1110
rect 155 830 165 1100
rect 185 830 245 1100
rect 265 830 275 1100
rect 155 820 275 830
rect 335 1100 375 1110
rect 335 830 345 1100
rect 365 830 375 1100
rect 335 820 375 830
rect 435 1100 555 1110
rect 435 830 445 1100
rect 465 830 525 1100
rect 545 830 555 1100
rect 435 820 555 830
rect 615 1100 655 1110
rect 615 830 625 1100
rect 645 830 655 1100
rect 615 820 655 830
rect 715 1100 835 1110
rect 715 830 725 1100
rect 745 830 805 1100
rect 825 830 835 1100
rect 715 820 835 830
rect 895 1100 935 1110
rect 895 830 905 1100
rect 925 830 935 1100
rect 895 820 935 830
rect 995 1100 1115 1110
rect 995 830 1005 1100
rect 1025 830 1085 1100
rect 1105 830 1115 1100
rect 995 820 1115 830
rect 1175 1100 1215 1110
rect 1175 830 1185 1100
rect 1205 830 1215 1100
rect 1175 820 1215 830
rect 1275 1100 1315 1110
rect 1275 830 1285 1100
rect 1305 830 1315 1100
rect 1275 820 1315 830
rect 65 800 85 820
rect 345 800 365 820
rect 625 800 645 820
rect 905 800 925 820
rect 1185 800 1205 820
rect 5 740 45 750
rect 5 720 15 740
rect 35 720 45 740
rect 5 710 45 720
rect 1225 740 1265 750
rect 1225 720 1235 740
rect 1255 720 1265 740
rect 1225 710 1265 720
rect 65 690 85 710
rect 345 690 365 700
rect 625 690 645 700
rect 905 690 925 700
rect 1185 690 1205 700
rect -45 680 -5 690
rect -45 410 -35 680
rect -15 410 -5 680
rect -45 400 -5 410
rect 55 680 95 690
rect 55 410 65 680
rect 85 410 95 680
rect 55 400 95 410
rect 155 680 195 690
rect 155 410 165 680
rect 185 410 195 680
rect 155 400 195 410
rect 235 680 275 690
rect 235 410 245 680
rect 265 410 275 680
rect 235 400 275 410
rect 335 680 375 690
rect 335 410 345 680
rect 365 410 375 680
rect 335 400 375 410
rect 435 680 475 690
rect 435 410 445 680
rect 465 410 475 680
rect 435 400 475 410
rect 515 680 555 690
rect 515 410 525 680
rect 545 410 555 680
rect 515 400 555 410
rect 615 680 655 690
rect 615 410 625 680
rect 645 410 655 680
rect 615 400 655 410
rect 715 680 755 690
rect 715 410 725 680
rect 745 410 755 680
rect 715 400 755 410
rect 795 680 835 690
rect 795 410 805 680
rect 825 410 835 680
rect 795 400 835 410
rect 895 680 935 690
rect 895 410 905 680
rect 925 410 935 680
rect 895 400 935 410
rect 995 680 1035 690
rect 995 410 1005 680
rect 1025 410 1035 680
rect 995 400 1035 410
rect 1075 680 1115 690
rect 1075 410 1085 680
rect 1105 410 1115 680
rect 1075 400 1115 410
rect 1175 680 1215 690
rect 1175 410 1185 680
rect 1205 410 1215 680
rect 1175 400 1215 410
rect 1275 680 1315 690
rect 1275 410 1285 680
rect 1305 410 1315 680
rect 1275 400 1315 410
rect 175 355 195 400
rect 175 345 215 355
rect 175 325 185 345
rect 205 325 215 345
rect 175 315 215 325
rect 245 335 265 400
rect 455 355 475 400
rect 455 345 515 355
rect 455 335 485 345
rect 245 325 485 335
rect 505 325 515 345
rect 245 315 515 325
rect 535 335 555 400
rect 615 345 655 355
rect 615 335 625 345
rect 535 325 625 335
rect 645 335 655 345
rect 725 335 745 400
rect 805 355 825 400
rect 645 325 745 335
rect 535 315 745 325
rect 765 345 825 355
rect 765 325 775 345
rect 795 335 825 345
rect 1005 335 1025 400
rect 1075 355 1095 400
rect 795 325 1025 335
rect 765 315 1025 325
rect 1055 345 1095 355
rect 1055 325 1065 345
rect 1085 325 1095 345
rect 1055 315 1095 325
rect 175 295 195 315
rect 245 295 265 315
rect 455 295 475 315
rect 535 295 555 315
rect 725 295 745 315
rect 805 295 825 315
rect 1005 295 1025 315
rect 1075 295 1095 315
rect -45 285 -5 295
rect -45 15 -35 285
rect -15 15 -5 285
rect -45 5 -5 15
rect 55 285 95 295
rect 55 15 65 285
rect 85 15 95 285
rect 55 5 95 15
rect 155 285 195 295
rect 155 15 165 285
rect 185 15 195 285
rect 155 5 195 15
rect 235 285 275 295
rect 235 15 245 285
rect 265 15 275 285
rect 235 5 275 15
rect 335 285 375 295
rect 335 15 345 285
rect 365 15 375 285
rect 335 5 375 15
rect 435 285 475 295
rect 435 15 445 285
rect 465 15 475 285
rect 435 5 475 15
rect 515 285 555 295
rect 515 15 525 285
rect 545 15 555 285
rect 515 5 555 15
rect 615 285 655 295
rect 615 15 625 285
rect 645 15 655 285
rect 615 5 655 15
rect 715 285 755 295
rect 715 15 725 285
rect 745 15 755 285
rect 715 5 755 15
rect 795 285 835 295
rect 795 15 805 285
rect 825 15 835 285
rect 795 5 835 15
rect 895 285 935 295
rect 895 15 905 285
rect 925 15 935 285
rect 895 5 935 15
rect 995 285 1035 295
rect 995 15 1005 285
rect 1025 15 1035 285
rect 995 5 1035 15
rect 1075 285 1115 295
rect 1075 15 1085 285
rect 1105 15 1115 285
rect 1075 5 1115 15
rect 1175 285 1215 295
rect 1175 15 1185 285
rect 1205 15 1215 285
rect 1175 5 1215 15
rect 1275 285 1315 295
rect 1275 15 1285 285
rect 1305 15 1315 285
rect 1275 5 1315 15
rect 5 -25 45 -15
rect 5 -45 15 -25
rect 35 -45 45 -25
rect 5 -55 45 -45
rect 65 -110 85 5
rect 345 -110 365 5
rect 625 -110 645 5
rect 905 -110 925 5
rect 1185 -110 1205 5
rect 1225 -25 1265 -15
rect 1225 -45 1235 -25
rect 1255 -45 1265 -25
rect 1225 -55 1265 -45
rect -45 -120 -5 -110
rect -45 -390 -35 -120
rect -15 -390 -5 -120
rect -45 -400 -5 -390
rect 55 -120 95 -110
rect 55 -390 65 -120
rect 85 -390 95 -120
rect 55 -400 95 -390
rect 155 -120 275 -110
rect 155 -390 165 -120
rect 185 -390 245 -120
rect 265 -390 275 -120
rect 155 -400 275 -390
rect 335 -120 375 -110
rect 335 -390 345 -120
rect 365 -390 375 -120
rect 335 -400 375 -390
rect 435 -120 555 -110
rect 435 -390 445 -120
rect 465 -390 525 -120
rect 545 -390 555 -120
rect 435 -400 555 -390
rect 615 -120 655 -110
rect 615 -390 625 -120
rect 645 -390 655 -120
rect 615 -400 655 -390
rect 715 -120 835 -110
rect 715 -390 725 -120
rect 745 -390 805 -120
rect 825 -390 835 -120
rect 715 -400 835 -390
rect 895 -120 935 -110
rect 895 -390 905 -120
rect 925 -390 935 -120
rect 895 -400 935 -390
rect 995 -120 1115 -110
rect 995 -390 1005 -120
rect 1025 -390 1085 -120
rect 1105 -390 1115 -120
rect 995 -400 1115 -390
rect 1175 -120 1215 -110
rect 1175 -390 1185 -120
rect 1205 -390 1215 -120
rect 1175 -400 1215 -390
rect 1275 -120 1315 -110
rect 1275 -390 1285 -120
rect 1305 -390 1315 -120
rect 1275 -400 1315 -390
rect 5 -430 45 -420
rect 5 -450 15 -430
rect 35 -450 45 -430
rect 5 -460 45 -450
rect 1225 -430 1265 -420
rect 1225 -450 1235 -430
rect 1255 -450 1265 -430
rect 1225 -460 1265 -450
<< viali >>
rect -35 1780 -15 2050
rect 165 1780 185 2050
rect 245 1780 265 2050
rect 445 1780 465 2050
rect 525 1780 545 2050
rect 725 1780 745 2050
rect 805 1780 825 2050
rect 1005 1780 1025 2050
rect 1085 1780 1105 2050
rect 1285 1780 1305 2050
rect -35 1310 -15 1580
rect 1285 1310 1305 1580
rect -35 830 -15 1100
rect 165 830 185 1100
rect 245 830 265 1100
rect 445 830 465 1100
rect 525 830 545 1100
rect 725 830 745 1100
rect 805 830 825 1100
rect 1005 830 1025 1100
rect 1085 830 1105 1100
rect 1285 830 1305 1100
rect 185 325 205 345
rect 625 325 645 345
rect 1065 325 1085 345
rect -35 -390 -15 -120
rect 165 -390 185 -120
rect 245 -390 265 -120
rect 445 -390 465 -120
rect 525 -390 545 -120
rect 725 -390 745 -120
rect 805 -390 825 -120
rect 1005 -390 1025 -120
rect 1085 -390 1105 -120
rect 1285 -390 1305 -120
<< metal1 >>
rect 175 345 1095 355
rect 175 325 185 345
rect 205 340 625 345
rect 205 325 215 340
rect 175 315 215 325
rect 615 325 625 340
rect 645 340 1065 345
rect 645 325 655 340
rect 615 315 655 325
rect 1055 325 1065 340
rect 1085 325 1095 345
rect 1055 315 1095 325
<< end >>
